module formal_bind;
    bind design_top.dut.irf formal_spec chk0 (.clk(CLK),
                                           .rst(1'b0),
                                           .reg0 ('b0),
                                           .reg1 (Q[1]),
                                           .reg2 (Q[2]),
                                           .reg3 (Q[3]),
                                           .reg4 (Q[4]),
                                           .reg5 (Q[5]),
                                           .reg6 (Q[6]),
                                           .reg7 (Q[7]),
                                           .reg8 (Q[8]),
                                           .reg9 (Q[9]),
                                           .reg10(Q[10]),
                                           .reg11(Q[11]),
                                           .reg12(Q[12]),
                                           .reg13(Q[13]),
                                           .reg14(Q[14]),
                                           .reg15(Q[15]),
                                           .reg16(Q[16]),
                                           .reg17(Q[17]),
                                           .reg18(Q[18]),
                                           .reg19(Q[19]),
                                           .reg20(Q[20]),
                                           .reg21(Q[21]),
                                           .reg22(Q[22]),
                                           .reg23(Q[23]),
                                           .reg24(Q[24]),
                                           .reg25(Q[25]),
                                           .reg26(Q[26]),
                                           .reg27(Q[27]),
                                           .reg28(Q[28]),
                                           .reg29(Q[29]),
                                           .reg30(Q[30]),
                                           .reg31(Q[31]));
endmodule
