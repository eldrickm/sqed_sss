module vscale_checker_bind;

    bind picorv32 picorv32_checker chk0 (.clk(clk),
                                         .rst(1'b0),
                                         .reg0 (cpuregs[0]),
                                         .reg1 (cpuregs[1]),
                                         .reg2 (cpuregs[2]),
                                         .reg3 (cpuregs[3]),
                                         .reg4 (cpuregs[4]),
                                         .reg5 (cpuregs[5]),
                                         .reg6 (cpuregs[6]),
                                         .reg7 (cpuregs[7]),
                                         .reg8 (cpuregs[8]),
                                         .reg9 (cpuregs[9]),
                                         .reg10(cpuregs[10]),
                                         .reg11(cpuregs[11]),
                                         .reg12(cpuregs[12]),
                                         .reg13(cpuregs[13]),
                                         .reg14(cpuregs[14]),
                                         .reg15(cpuregs[15]),
                                         .reg16(cpuregs[16]),
                                         .reg17(cpuregs[17]),
                                         .reg18(cpuregs[18]),
                                         .reg19(cpuregs[19]),
                                         .reg20(cpuregs[20]),
                                         .reg21(cpuregs[21]),
                                         .reg22(cpuregs[22]),
                                         .reg23(cpuregs[23]),
                                         .reg24(cpuregs[24]),
                                         .reg25(cpuregs[25]),
                                         .reg26(cpuregs[26]),
                                         .reg27(cpuregs[27]),
                                         .reg28(cpuregs[28]),
                                         .reg29(cpuregs[29]),
                                         .reg30(cpuregs[30]),
                                         .reg31(cpuregs[31]));

endmodule
