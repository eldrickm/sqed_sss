module Queue_5_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 34016:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 34017:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 34018:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input  [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input  [7:0]  io_enq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [7:0]  io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output        io_deq_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output        io_deq_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg [7:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [7:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [7:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg  ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34022:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34023:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 34024:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 34025:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 34026:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 34027:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 34028:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 34029:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 34032:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 34047:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 34053:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 34056:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_param_MPORT_data = 2'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_sink_MPORT_data = 1'h0;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_denied_MPORT_data = 1'h0;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 34062:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 34060:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34072:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34071:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34070:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34069:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34068:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34067:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34066:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34065:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34022:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34022:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 34035:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 34048:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34023:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34023:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 34050:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 34054:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 34024:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 34024:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 34057:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 34058:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 39472:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 39473:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 39474:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [31:0] io_enq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output        io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [31:0] io_deq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39478:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39479:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39480:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 39481:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 39482:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 39483:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 39484:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 39485:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 39488:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 39503:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 39509:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 39512:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_param_MPORT_data = 3'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_source_MPORT_data = 1'h0;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 39518:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 39516:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39528:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39527:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39526:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39525:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39524:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39523:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39522:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39521:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39478:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39478:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 39491:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 39504:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39479:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39479:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 39506:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 39510:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39480:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39480:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 39513:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 39514:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_7_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 39536:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 39537:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 39538:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [1:0]  io_enq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_enq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [2:0]  io_enq_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_enq_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output        io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [2:0]  io_deq_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output        io_deq_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg [2:0] ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [2:0] ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [2:0] ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39542:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39543:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39544:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 39545:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 39546:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 39547:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 39548:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 39549:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 39552:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 39567:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 39573:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 39576:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_sink_MPORT_data = io_enq_bits_sink;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 39582:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 39580:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39592:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39591:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39590:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39589:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39588:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39587:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39586:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39585:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39542:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39542:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 39555:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 39568:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39543:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39543:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 39570:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 39574:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39544:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39544:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 39577:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 39578:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HellaPeekingArbiter_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 369278:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 369279:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 369280:4]
  output        io_in_1_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input         io_in_1_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [2:0]  io_in_1_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [2:0]  io_in_1_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [3:0]  io_in_1_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [3:0]  io_in_1_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [63:0] io_in_1_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input         io_in_1_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [7:0]  io_in_1_bits_union, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input         io_in_1_bits_last, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output        io_in_4_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input         io_in_4_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [2:0]  io_in_4_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [2:0]  io_in_4_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [3:0]  io_in_4_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [3:0]  io_in_4_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [31:0] io_in_4_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [63:0] io_in_4_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input         io_in_4_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input  [7:0]  io_in_4_bits_union, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input         io_in_4_bits_last, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  input         io_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output        io_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output [2:0]  io_out_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output [3:0]  io_out_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output [3:0]  io_out_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output [31:0] io_out_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output [63:0] io_out_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output        io_out_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output [7:0]  io_out_bits_union, // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
  output        io_out_bits_last // @[chipyard.TestHarness.SmallBoomConfig.fir 369281:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockIdx; // @[Arbiters.scala 25:20 chipyard.TestHarness.SmallBoomConfig.fir 369286:4]
  reg  locked; // @[Arbiters.scala 26:19 chipyard.TestHarness.SmallBoomConfig.fir 369287:4]
  wire [2:0] choice = io_in_1_valid ? 3'h1 : 3'h4; // @[Mux.scala 47:69 chipyard.TestHarness.SmallBoomConfig.fir 369290:4]
  wire [2:0] chosen = locked ? lockIdx : choice; // @[Arbiters.scala 36:19 chipyard.TestHarness.SmallBoomConfig.fir 369292:4]
  wire  _io_in_1_ready_T = chosen == 3'h1; // @[Arbiters.scala 39:46 chipyard.TestHarness.SmallBoomConfig.fir 369296:4]
  wire  _io_in_4_ready_T = chosen == 3'h4; // @[Arbiters.scala 39:46 chipyard.TestHarness.SmallBoomConfig.fir 369305:4]
  wire [2:0] _GEN_14 = 3'h1 == chosen ? 3'h3 : 3'h4; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [2:0] _GEN_15 = 3'h1 == chosen ? io_in_1_bits_opcode : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [2:0] _GEN_16 = 3'h1 == chosen ? io_in_1_bits_param : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [3:0] _GEN_17 = 3'h1 == chosen ? io_in_1_bits_size : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [3:0] _GEN_18 = 3'h1 == chosen ? io_in_1_bits_source : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [63:0] _GEN_20 = 3'h1 == chosen ? io_in_1_bits_data : 64'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [7:0] _GEN_22 = 3'h1 == chosen ? io_in_1_bits_union : 8'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire  _GEN_23 = 3'h1 == chosen ? io_in_1_bits_last : 1'h1; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire  _GEN_25 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_valid; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [2:0] _GEN_26 = 3'h2 == chosen ? 3'h2 : _GEN_14; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [2:0] _GEN_27 = 3'h2 == chosen ? 3'h0 : _GEN_15; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [2:0] _GEN_28 = 3'h2 == chosen ? 3'h0 : _GEN_16; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [3:0] _GEN_29 = 3'h2 == chosen ? 4'h0 : _GEN_17; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [3:0] _GEN_30 = 3'h2 == chosen ? 4'h0 : _GEN_18; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [63:0] _GEN_32 = 3'h2 == chosen ? 64'h0 : _GEN_20; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire  _GEN_33 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_bits_corrupt; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [7:0] _GEN_34 = 3'h2 == chosen ? 8'h0 : _GEN_22; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire  _GEN_37 = 3'h3 == chosen ? 1'h0 : _GEN_25; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [2:0] _GEN_38 = 3'h3 == chosen ? 3'h1 : _GEN_26; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [2:0] _GEN_39 = 3'h3 == chosen ? 3'h0 : _GEN_27; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [2:0] _GEN_40 = 3'h3 == chosen ? 3'h0 : _GEN_28; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [3:0] _GEN_41 = 3'h3 == chosen ? 4'h0 : _GEN_29; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [3:0] _GEN_42 = 3'h3 == chosen ? 4'h0 : _GEN_30; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [63:0] _GEN_44 = 3'h3 == chosen ? 64'h0 : _GEN_32; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire  _GEN_45 = 3'h3 == chosen ? 1'h0 : _GEN_33; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire [7:0] _GEN_46 = 3'h3 == chosen ? 8'h0 : _GEN_34; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369310:4]
  wire  _T_1 = ~locked; // @[Arbiters.scala 59:11 chipyard.TestHarness.SmallBoomConfig.fir 369312:6]
  wire  _GEN_61 = _T_1 | locked; // @[Arbiters.scala 59:50 chipyard.TestHarness.SmallBoomConfig.fir 369314:6 Arbiters.scala 61:14 chipyard.TestHarness.SmallBoomConfig.fir 369316:8 Arbiters.scala 26:19 chipyard.TestHarness.SmallBoomConfig.fir 369287:4]
  assign io_in_1_ready = io_out_ready & _io_in_1_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.SmallBoomConfig.fir 369297:4]
  assign io_in_4_ready = io_out_ready & _io_in_4_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.SmallBoomConfig.fir 369306:4]
  assign io_out_valid = 3'h4 == chosen ? io_in_4_valid : _GEN_37; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_chanId = 3'h4 == chosen ? 3'h0 : _GEN_38; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_opcode = 3'h4 == chosen ? io_in_4_bits_opcode : _GEN_39; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_param = 3'h4 == chosen ? io_in_4_bits_param : _GEN_40; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_size = 3'h4 == chosen ? io_in_4_bits_size : _GEN_41; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_source = 3'h4 == chosen ? io_in_4_bits_source : _GEN_42; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_address = 3'h4 == chosen ? io_in_4_bits_address : 32'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_data = 3'h4 == chosen ? io_in_4_bits_data : _GEN_44; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_corrupt = 3'h4 == chosen ? io_in_4_bits_corrupt : _GEN_45; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_union = 3'h4 == chosen ? io_in_4_bits_union : _GEN_46; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  assign io_out_bits_last = 3'h4 == chosen ? io_in_4_bits_last : 3'h3 == chosen | (3'h2 == chosen | _GEN_23); // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369308:4]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiters.scala 25:20 chipyard.TestHarness.SmallBoomConfig.fir 369286:4]
      lockIdx <= 3'h0; // @[Arbiters.scala 25:20 chipyard.TestHarness.SmallBoomConfig.fir 369286:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.SmallBoomConfig.fir 369311:4]
      if (_T_1) begin // @[Arbiters.scala 59:50 chipyard.TestHarness.SmallBoomConfig.fir 369314:6]
        if (io_in_1_valid) begin // @[Mux.scala 47:69 chipyard.TestHarness.SmallBoomConfig.fir 369290:4]
          lockIdx <= 3'h1;
        end else begin
          lockIdx <= 3'h4;
        end
      end
    end
    if (reset) begin // @[Arbiters.scala 26:19 chipyard.TestHarness.SmallBoomConfig.fir 369287:4]
      locked <= 1'h0; // @[Arbiters.scala 26:19 chipyard.TestHarness.SmallBoomConfig.fir 369287:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.SmallBoomConfig.fir 369311:4]
      if (io_out_bits_last) begin // @[Arbiters.scala 64:35 chipyard.TestHarness.SmallBoomConfig.fir 369318:6]
        locked <= 1'h0; // @[Arbiters.scala 65:14 chipyard.TestHarness.SmallBoomConfig.fir 369319:8]
      end else begin
        locked <= _GEN_61;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockIdx = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  locked = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericSerializer_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 369323:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 369324:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 369325:4]
  output        io_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input         io_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input  [2:0]  io_in_bits_chanId, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input  [2:0]  io_in_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input  [2:0]  io_in_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input  [3:0]  io_in_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input  [3:0]  io_in_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input  [31:0] io_in_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input  [63:0] io_in_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input         io_in_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input  [7:0]  io_in_bits_union, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input         io_in_bits_last, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  input         io_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  output        io_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
  output [3:0]  io_out_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 369326:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [122:0] data; // @[Serdes.scala 175:17 chipyard.TestHarness.SmallBoomConfig.fir 369328:4]
  reg  sending; // @[Serdes.scala 177:24 chipyard.TestHarness.SmallBoomConfig.fir 369329:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369330:4]
  reg [4:0] sendCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369331:4]
  wire  wrap_wrap = sendCount == 5'h1e; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 369335:6]
  wire [4:0] _wrap_value_T_1 = sendCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 369337:6]
  wire  sendDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 369334:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 369342:6 chipyard.TestHarness.SmallBoomConfig.fir 369333:4]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369349:4]
  wire [122:0] _data_T = {io_in_bits_chanId,io_in_bits_opcode,io_in_bits_param,io_in_bits_size,io_in_bits_source,
    io_in_bits_address,io_in_bits_data,io_in_bits_corrupt,io_in_bits_union,io_in_bits_last}; // @[Serdes.scala 185:24 chipyard.TestHarness.SmallBoomConfig.fir 369359:6]
  wire  _GEN_4 = _T_1 | sending; // @[Serdes.scala 184:23 chipyard.TestHarness.SmallBoomConfig.fir 369350:4 Serdes.scala 186:13 chipyard.TestHarness.SmallBoomConfig.fir 369361:6 Serdes.scala 177:24 chipyard.TestHarness.SmallBoomConfig.fir 369329:4]
  wire [122:0] _data_T_1 = {{4'd0}, data[122:4]}; // @[Serdes.scala 189:39 chipyard.TestHarness.SmallBoomConfig.fir 369365:6]
  assign io_in_ready = ~sending; // @[Serdes.scala 180:18 chipyard.TestHarness.SmallBoomConfig.fir 369344:4]
  assign io_out_valid = sending; // @[Serdes.scala 181:16 chipyard.TestHarness.SmallBoomConfig.fir 369346:4]
  assign io_out_bits = data[3:0]; // @[Serdes.scala 182:22 chipyard.TestHarness.SmallBoomConfig.fir 369347:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 189:24 chipyard.TestHarness.SmallBoomConfig.fir 369364:4]
      data <= _data_T_1; // @[Serdes.scala 189:31 chipyard.TestHarness.SmallBoomConfig.fir 369366:6]
    end else if (_T_1) begin // @[Serdes.scala 184:23 chipyard.TestHarness.SmallBoomConfig.fir 369350:4]
      data <= _data_T; // @[Serdes.scala 185:10 chipyard.TestHarness.SmallBoomConfig.fir 369360:6]
    end
    if (reset) begin // @[Serdes.scala 177:24 chipyard.TestHarness.SmallBoomConfig.fir 369329:4]
      sending <= 1'h0; // @[Serdes.scala 177:24 chipyard.TestHarness.SmallBoomConfig.fir 369329:4]
    end else if (sendDone) begin // @[Serdes.scala 191:19 chipyard.TestHarness.SmallBoomConfig.fir 369368:4]
      sending <= 1'h0; // @[Serdes.scala 191:29 chipyard.TestHarness.SmallBoomConfig.fir 369369:6]
    end else begin
      sending <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369331:4]
      sendCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369331:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 369334:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.SmallBoomConfig.fir 369339:6]
        sendCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.SmallBoomConfig.fir 369340:8]
      end else begin
        sendCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 369338:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data = _RAND_0[122:0];
  _RAND_1 = {1{`RANDOM}};
  sending = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sendCount = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericDeserializer_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 369372:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 369373:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 369374:4]
  output        io_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  input         io_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  input  [3:0]  io_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  input         io_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output        io_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output [2:0]  io_out_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output [3:0]  io_out_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output [3:0]  io_out_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output [31:0] io_out_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output [63:0] io_out_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output        io_out_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
  output [7:0]  io_out_bits_union // @[chipyard.TestHarness.SmallBoomConfig.fir 369375:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] data_0; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_1; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_2; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_3; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_4; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_5; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_6; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_7; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_8; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_9; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_10; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_11; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_12; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_13; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_14; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_15; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_16; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_17; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_18; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_19; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_20; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_21; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_22; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_23; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_24; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_25; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_26; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_27; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_28; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_29; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg [3:0] data_30; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369377:4]
  reg  receiving; // @[Serdes.scala 204:26 chipyard.TestHarness.SmallBoomConfig.fir 369378:4]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369379:4]
  reg [4:0] recvCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369380:4]
  wire  wrap_wrap = recvCount == 5'h1e; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 369384:6]
  wire [4:0] _wrap_value_T_1 = recvCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 369386:6]
  wire  recvDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 369383:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 369391:6 chipyard.TestHarness.SmallBoomConfig.fir 369382:4]
  wire [27:0] io_out_bits_lo_lo = {data_6,data_5,data_4,data_3,data_2,data_1,data_0}; // @[Serdes.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 369401:4]
  wire [59:0] io_out_bits_lo = {data_14,data_13,data_12,data_11,data_10,data_9,data_8,data_7,io_out_bits_lo_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 369409:4]
  wire [31:0] io_out_bits_hi_lo = {data_22,data_21,data_20,data_19,data_18,data_17,data_16,data_15}; // @[Serdes.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 369416:4]
  wire [123:0] _io_out_bits_T = {data_30,data_29,data_28,data_27,data_26,data_25,data_24,data_23,io_out_bits_hi_lo,
    io_out_bits_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 369425:4]
  wire  _GEN_65 = recvDone ? 1'h0 : receiving; // @[Serdes.scala 215:19 chipyard.TestHarness.SmallBoomConfig.fir 369463:4 Serdes.scala 215:31 chipyard.TestHarness.SmallBoomConfig.fir 369464:6 Serdes.scala 204:26 chipyard.TestHarness.SmallBoomConfig.fir 369378:4]
  wire  _T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369466:4]
  wire  _GEN_66 = _T_2 | _GEN_65; // @[Serdes.scala 217:24 chipyard.TestHarness.SmallBoomConfig.fir 369467:4 Serdes.scala 217:36 chipyard.TestHarness.SmallBoomConfig.fir 369468:6]
  assign io_in_ready = receiving; // @[Serdes.scala 207:15 chipyard.TestHarness.SmallBoomConfig.fir 369393:4]
  assign io_out_valid = ~receiving; // @[Serdes.scala 208:19 chipyard.TestHarness.SmallBoomConfig.fir 369394:4]
  assign io_out_bits_chanId = _io_out_bits_T[122:120]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369447:4]
  assign io_out_bits_opcode = _io_out_bits_T[119:117]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369445:4]
  assign io_out_bits_param = _io_out_bits_T[116:114]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369443:4]
  assign io_out_bits_size = _io_out_bits_T[113:110]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369441:4]
  assign io_out_bits_source = _io_out_bits_T[109:106]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369439:4]
  assign io_out_bits_address = _io_out_bits_T[105:74]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369437:4]
  assign io_out_bits_data = _io_out_bits_T[73:10]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369435:4]
  assign io_out_bits_corrupt = _io_out_bits_T[9]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369433:4]
  assign io_out_bits_union = _io_out_bits_T[8:1]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369431:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h0 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_0 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h1 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_1 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h2 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_2 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h3 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_3 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h4 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_4 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h5 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_5 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h6 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_6 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h7 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_7 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h8 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_8 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h9 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_9 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'ha == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_10 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'hb == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_11 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'hc == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_12 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'hd == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_13 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'he == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_14 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'hf == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_15 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h10 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_16 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h11 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_17 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h12 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_18 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h13 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_19 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h14 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_20 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h15 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_21 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h16 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_22 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h17 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_23 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h18 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_24 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h19 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_25 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h1a == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_26 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h1b == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_27 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h1c == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_28 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h1d == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_29 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369460:4]
      if (5'h1e == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
        data_30 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369461:6]
      end
    end
    receiving <= reset | _GEN_66; // @[Serdes.scala 204:26 chipyard.TestHarness.SmallBoomConfig.fir 369378:4 Serdes.scala 204:26 chipyard.TestHarness.SmallBoomConfig.fir 369378:4]
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369380:4]
      recvCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369380:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 369383:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.SmallBoomConfig.fir 369388:6]
        recvCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.SmallBoomConfig.fir 369389:8]
      end else begin
        recvCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 369387:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  data_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  data_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  data_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  data_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  data_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  data_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  data_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  data_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  data_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  data_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  data_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  data_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  data_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  data_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  data_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  data_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  data_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  data_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  data_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  data_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  data_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  data_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  data_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  data_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  data_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  data_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  data_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  data_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  data_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  data_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  receiving = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  recvCount = _RAND_32[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SerialAdapter_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 380448:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 380449:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 380450:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  output [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  output [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 380451:4]
  output        io_serial_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 380452:4]
  input         io_serial_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 380452:4]
  input  [31:0] io_serial_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 380452:4]
  input         io_serial_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 380452:4]
  output        io_serial_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 380452:4]
  output [31:0] io_serial_out_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 380452:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cmd; // @[SerialAdapter.scala 86:16 chipyard.TestHarness.SmallBoomConfig.fir 380461:4]
  reg [63:0] addr; // @[SerialAdapter.scala 87:17 chipyard.TestHarness.SmallBoomConfig.fir 380462:4]
  reg [63:0] len; // @[SerialAdapter.scala 88:16 chipyard.TestHarness.SmallBoomConfig.fir 380463:4]
  reg [31:0] body_0; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.SmallBoomConfig.fir 380464:4]
  reg [31:0] body_1; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.SmallBoomConfig.fir 380464:4]
  reg [1:0] bodyValid; // @[SerialAdapter.scala 90:22 chipyard.TestHarness.SmallBoomConfig.fir 380465:4]
  reg  idx; // @[SerialAdapter.scala 91:16 chipyard.TestHarness.SmallBoomConfig.fir 380466:4]
  reg [3:0] state; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.SmallBoomConfig.fir 380467:4]
  wire  _io_serial_in_ready_T = state == 4'h0; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380468:4]
  wire  _io_serial_in_ready_T_1 = state == 4'h1; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380469:4]
  wire  _io_serial_in_ready_T_2 = state == 4'h2; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380470:4]
  wire  _io_serial_in_ready_T_3 = state == 4'h6; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380471:4]
  wire  _io_serial_in_ready_T_4 = _io_serial_in_ready_T | _io_serial_in_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380472:4]
  wire  _io_serial_in_ready_T_5 = _io_serial_in_ready_T_4 | _io_serial_in_ready_T_2; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380473:4]
  wire  _io_serial_out_valid_T = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.SmallBoomConfig.fir 380476:4]
  wire [28:0] beatAddr = addr[31:3]; // @[SerialAdapter.scala 103:22 chipyard.TestHarness.SmallBoomConfig.fir 380479:4]
  wire [28:0] nextAddr_hi = beatAddr + 29'h1; // @[SerialAdapter.scala 104:31 chipyard.TestHarness.SmallBoomConfig.fir 380481:4]
  wire [31:0] nextAddr = {nextAddr_hi,3'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380482:4]
  wire [3:0] wmask_lo = bodyValid[0] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.SmallBoomConfig.fir 380486:4]
  wire [3:0] wmask_hi = bodyValid[1] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.SmallBoomConfig.fir 380488:4]
  wire [7:0] wmask = {wmask_hi,wmask_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380489:4]
  wire [63:0] _GEN_55 = {{32'd0}, nextAddr}; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.SmallBoomConfig.fir 380490:4]
  wire [63:0] addr_size = _GEN_55 - addr; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.SmallBoomConfig.fir 380491:4]
  wire [63:0] len_size_hi = len + 64'h1; // @[SerialAdapter.scala 108:26 chipyard.TestHarness.SmallBoomConfig.fir 380493:4]
  wire [65:0] len_size = {len_size_hi,2'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380494:4]
  wire [65:0] _GEN_56 = {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 380495:4]
  wire  _raw_size_T = len_size < _GEN_56; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 380495:4]
  wire [65:0] raw_size = _raw_size_T ? len_size : {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:21 chipyard.TestHarness.SmallBoomConfig.fir 380496:4]
  wire  _rsize_T = 66'h1 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 380497:4]
  wire [1:0] _rsize_T_1 = _rsize_T ? 2'h0 : 2'h3; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 380498:4]
  wire  _rsize_T_2 = 66'h2 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 380499:4]
  wire [1:0] _rsize_T_3 = _rsize_T_2 ? 2'h1 : _rsize_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 380500:4]
  wire  _rsize_T_4 = 66'h4 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 380501:4]
  wire [1:0] rsize = _rsize_T_4 ? 2'h2 : _rsize_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 380502:4]
  wire [1:0] _pow2size_T_66 = raw_size[0] + raw_size[1]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380569:4]
  wire [1:0] _pow2size_T_68 = raw_size[2] + raw_size[3]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380571:4]
  wire [2:0] _pow2size_T_70 = _pow2size_T_66 + _pow2size_T_68; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380573:4]
  wire [1:0] _pow2size_T_72 = raw_size[4] + raw_size[5]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380575:4]
  wire [1:0] _pow2size_T_74 = raw_size[6] + raw_size[7]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380577:4]
  wire [2:0] _pow2size_T_76 = _pow2size_T_72 + _pow2size_T_74; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380579:4]
  wire [3:0] _pow2size_T_78 = _pow2size_T_70 + _pow2size_T_76; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380581:4]
  wire [1:0] _pow2size_T_80 = raw_size[8] + raw_size[9]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380583:4]
  wire [1:0] _pow2size_T_82 = raw_size[10] + raw_size[11]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380585:4]
  wire [2:0] _pow2size_T_84 = _pow2size_T_80 + _pow2size_T_82; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380587:4]
  wire [1:0] _pow2size_T_86 = raw_size[12] + raw_size[13]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380589:4]
  wire [1:0] _pow2size_T_88 = raw_size[14] + raw_size[15]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380591:4]
  wire [2:0] _pow2size_T_90 = _pow2size_T_86 + _pow2size_T_88; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380593:4]
  wire [3:0] _pow2size_T_92 = _pow2size_T_84 + _pow2size_T_90; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380595:4]
  wire [4:0] _pow2size_T_94 = _pow2size_T_78 + _pow2size_T_92; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380597:4]
  wire [1:0] _pow2size_T_96 = raw_size[16] + raw_size[17]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380599:4]
  wire [1:0] _pow2size_T_98 = raw_size[18] + raw_size[19]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380601:4]
  wire [2:0] _pow2size_T_100 = _pow2size_T_96 + _pow2size_T_98; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380603:4]
  wire [1:0] _pow2size_T_102 = raw_size[20] + raw_size[21]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380605:4]
  wire [1:0] _pow2size_T_104 = raw_size[22] + raw_size[23]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380607:4]
  wire [2:0] _pow2size_T_106 = _pow2size_T_102 + _pow2size_T_104; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380609:4]
  wire [3:0] _pow2size_T_108 = _pow2size_T_100 + _pow2size_T_106; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380611:4]
  wire [1:0] _pow2size_T_110 = raw_size[24] + raw_size[25]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380613:4]
  wire [1:0] _pow2size_T_112 = raw_size[26] + raw_size[27]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380615:4]
  wire [2:0] _pow2size_T_114 = _pow2size_T_110 + _pow2size_T_112; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380617:4]
  wire [1:0] _pow2size_T_116 = raw_size[28] + raw_size[29]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380619:4]
  wire [1:0] _pow2size_T_118 = raw_size[31] + raw_size[32]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380621:4]
  wire [1:0] _GEN_57 = {{1'd0}, raw_size[30]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380623:4]
  wire [2:0] _pow2size_T_120 = _GEN_57 + _pow2size_T_118; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380623:4]
  wire [2:0] _pow2size_T_122 = _pow2size_T_116 + _pow2size_T_120[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380625:4]
  wire [3:0] _pow2size_T_124 = _pow2size_T_114 + _pow2size_T_122; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380627:4]
  wire [4:0] _pow2size_T_126 = _pow2size_T_108 + _pow2size_T_124; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380629:4]
  wire [5:0] _pow2size_T_128 = _pow2size_T_94 + _pow2size_T_126; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380631:4]
  wire [1:0] _pow2size_T_130 = raw_size[33] + raw_size[34]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380633:4]
  wire [1:0] _pow2size_T_132 = raw_size[35] + raw_size[36]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380635:4]
  wire [2:0] _pow2size_T_134 = _pow2size_T_130 + _pow2size_T_132; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380637:4]
  wire [1:0] _pow2size_T_136 = raw_size[37] + raw_size[38]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380639:4]
  wire [1:0] _pow2size_T_138 = raw_size[39] + raw_size[40]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380641:4]
  wire [2:0] _pow2size_T_140 = _pow2size_T_136 + _pow2size_T_138; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380643:4]
  wire [3:0] _pow2size_T_142 = _pow2size_T_134 + _pow2size_T_140; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380645:4]
  wire [1:0] _pow2size_T_144 = raw_size[41] + raw_size[42]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380647:4]
  wire [1:0] _pow2size_T_146 = raw_size[43] + raw_size[44]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380649:4]
  wire [2:0] _pow2size_T_148 = _pow2size_T_144 + _pow2size_T_146; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380651:4]
  wire [1:0] _pow2size_T_150 = raw_size[45] + raw_size[46]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380653:4]
  wire [1:0] _pow2size_T_152 = raw_size[47] + raw_size[48]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380655:4]
  wire [2:0] _pow2size_T_154 = _pow2size_T_150 + _pow2size_T_152; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380657:4]
  wire [3:0] _pow2size_T_156 = _pow2size_T_148 + _pow2size_T_154; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380659:4]
  wire [4:0] _pow2size_T_158 = _pow2size_T_142 + _pow2size_T_156; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380661:4]
  wire [1:0] _pow2size_T_160 = raw_size[49] + raw_size[50]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380663:4]
  wire [1:0] _pow2size_T_162 = raw_size[51] + raw_size[52]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380665:4]
  wire [2:0] _pow2size_T_164 = _pow2size_T_160 + _pow2size_T_162; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380667:4]
  wire [1:0] _pow2size_T_166 = raw_size[53] + raw_size[54]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380669:4]
  wire [1:0] _pow2size_T_168 = raw_size[55] + raw_size[56]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380671:4]
  wire [2:0] _pow2size_T_170 = _pow2size_T_166 + _pow2size_T_168; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380673:4]
  wire [3:0] _pow2size_T_172 = _pow2size_T_164 + _pow2size_T_170; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380675:4]
  wire [1:0] _pow2size_T_174 = raw_size[57] + raw_size[58]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380677:4]
  wire [1:0] _pow2size_T_176 = raw_size[59] + raw_size[60]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380679:4]
  wire [2:0] _pow2size_T_178 = _pow2size_T_174 + _pow2size_T_176; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380681:4]
  wire [1:0] _pow2size_T_180 = raw_size[61] + raw_size[62]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380683:4]
  wire [1:0] _pow2size_T_182 = raw_size[64] + raw_size[65]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380685:4]
  wire [1:0] _GEN_58 = {{1'd0}, raw_size[63]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380687:4]
  wire [2:0] _pow2size_T_184 = _GEN_58 + _pow2size_T_182; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380687:4]
  wire [2:0] _pow2size_T_186 = _pow2size_T_180 + _pow2size_T_184[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380689:4]
  wire [3:0] _pow2size_T_188 = _pow2size_T_178 + _pow2size_T_186; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380691:4]
  wire [4:0] _pow2size_T_190 = _pow2size_T_172 + _pow2size_T_188; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380693:4]
  wire [5:0] _pow2size_T_192 = _pow2size_T_158 + _pow2size_T_190; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380695:4]
  wire [6:0] _pow2size_T_194 = _pow2size_T_128 + _pow2size_T_192; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380697:4]
  wire  pow2size = _pow2size_T_194 == 7'h1; // @[SerialAdapter.scala 113:37 chipyard.TestHarness.SmallBoomConfig.fir 380699:4]
  wire [2:0] byteAddr = pow2size ? addr[2:0] : 3'h0; // @[SerialAdapter.scala 114:21 chipyard.TestHarness.SmallBoomConfig.fir 380701:4]
  wire [31:0] put_acquire_address = {beatAddr, 3'h0}; // @[SerialAdapter.scala 117:19 chipyard.TestHarness.SmallBoomConfig.fir 380702:4]
  wire [63:0] put_acquire_data = {body_1,body_0}; // @[SerialAdapter.scala 118:10 chipyard.TestHarness.SmallBoomConfig.fir 380703:4]
  wire [31:0] get_acquire_address = {beatAddr,byteAddr}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380768:4]
  wire [2:0] _get_acquire_a_mask_sizeOH_T = {{1'd0}, rsize}; // @[Misc.scala 201:34 chipyard.TestHarness.SmallBoomConfig.fir 380834:4]
  wire [1:0] get_acquire_a_mask_sizeOH_shiftAmount = _get_acquire_a_mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 380835:4]
  wire [3:0] _get_acquire_a_mask_sizeOH_T_1 = 4'h1 << get_acquire_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 380836:4]
  wire [2:0] get_acquire_a_mask_sizeOH = _get_acquire_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 380838:4]
  wire  _get_acquire_a_mask_T = rsize >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 380839:4]
  wire  get_acquire_a_mask_size = get_acquire_a_mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 380840:4]
  wire  get_acquire_a_mask_bit = get_acquire_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 380841:4]
  wire  get_acquire_a_mask_nbit = ~get_acquire_a_mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 380842:4]
  wire  _get_acquire_a_mask_acc_T = get_acquire_a_mask_size & get_acquire_a_mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380844:4]
  wire  get_acquire_a_mask_acc = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380845:4]
  wire  _get_acquire_a_mask_acc_T_1 = get_acquire_a_mask_size & get_acquire_a_mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380847:4]
  wire  get_acquire_a_mask_acc_1 = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380848:4]
  wire  get_acquire_a_mask_size_1 = get_acquire_a_mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 380849:4]
  wire  get_acquire_a_mask_bit_1 = get_acquire_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 380850:4]
  wire  get_acquire_a_mask_nbit_1 = ~get_acquire_a_mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 380851:4]
  wire  get_acquire_a_mask_eq_2 = get_acquire_a_mask_nbit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380852:4]
  wire  _get_acquire_a_mask_acc_T_2 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380853:4]
  wire  get_acquire_a_mask_acc_2 = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380854:4]
  wire  get_acquire_a_mask_eq_3 = get_acquire_a_mask_nbit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380855:4]
  wire  _get_acquire_a_mask_acc_T_3 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380856:4]
  wire  get_acquire_a_mask_acc_3 = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380857:4]
  wire  get_acquire_a_mask_eq_4 = get_acquire_a_mask_bit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380858:4]
  wire  _get_acquire_a_mask_acc_T_4 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380859:4]
  wire  get_acquire_a_mask_acc_4 = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380860:4]
  wire  get_acquire_a_mask_eq_5 = get_acquire_a_mask_bit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380861:4]
  wire  _get_acquire_a_mask_acc_T_5 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380862:4]
  wire  get_acquire_a_mask_acc_5 = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380863:4]
  wire  get_acquire_a_mask_size_2 = get_acquire_a_mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 380864:4]
  wire  get_acquire_a_mask_bit_2 = get_acquire_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 380865:4]
  wire  get_acquire_a_mask_nbit_2 = ~get_acquire_a_mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 380866:4]
  wire  get_acquire_a_mask_eq_6 = get_acquire_a_mask_eq_2 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380867:4]
  wire  _get_acquire_a_mask_acc_T_6 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380868:4]
  wire  get_acquire_a_mask_lo_lo_lo = get_acquire_a_mask_acc_2 | _get_acquire_a_mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380869:4]
  wire  get_acquire_a_mask_eq_7 = get_acquire_a_mask_eq_2 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380870:4]
  wire  _get_acquire_a_mask_acc_T_7 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380871:4]
  wire  get_acquire_a_mask_lo_lo_hi = get_acquire_a_mask_acc_2 | _get_acquire_a_mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380872:4]
  wire  get_acquire_a_mask_eq_8 = get_acquire_a_mask_eq_3 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380873:4]
  wire  _get_acquire_a_mask_acc_T_8 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380874:4]
  wire  get_acquire_a_mask_lo_hi_lo = get_acquire_a_mask_acc_3 | _get_acquire_a_mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380875:4]
  wire  get_acquire_a_mask_eq_9 = get_acquire_a_mask_eq_3 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380876:4]
  wire  _get_acquire_a_mask_acc_T_9 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380877:4]
  wire  get_acquire_a_mask_lo_hi_hi = get_acquire_a_mask_acc_3 | _get_acquire_a_mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380878:4]
  wire  get_acquire_a_mask_eq_10 = get_acquire_a_mask_eq_4 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380879:4]
  wire  _get_acquire_a_mask_acc_T_10 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380880:4]
  wire  get_acquire_a_mask_hi_lo_lo = get_acquire_a_mask_acc_4 | _get_acquire_a_mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380881:4]
  wire  get_acquire_a_mask_eq_11 = get_acquire_a_mask_eq_4 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380882:4]
  wire  _get_acquire_a_mask_acc_T_11 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380883:4]
  wire  get_acquire_a_mask_hi_lo_hi = get_acquire_a_mask_acc_4 | _get_acquire_a_mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380884:4]
  wire  get_acquire_a_mask_eq_12 = get_acquire_a_mask_eq_5 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380885:4]
  wire  _get_acquire_a_mask_acc_T_12 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380886:4]
  wire  get_acquire_a_mask_hi_hi_lo = get_acquire_a_mask_acc_5 | _get_acquire_a_mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380887:4]
  wire  get_acquire_a_mask_eq_13 = get_acquire_a_mask_eq_5 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380888:4]
  wire  _get_acquire_a_mask_acc_T_13 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380889:4]
  wire  get_acquire_a_mask_hi_hi_hi = get_acquire_a_mask_acc_5 | _get_acquire_a_mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380890:4]
  wire [7:0] get_acquire_mask = {get_acquire_a_mask_hi_hi_hi,get_acquire_a_mask_hi_hi_lo,get_acquire_a_mask_hi_lo_hi,
    get_acquire_a_mask_hi_lo_lo,get_acquire_a_mask_lo_hi_hi,get_acquire_a_mask_lo_hi_lo,get_acquire_a_mask_lo_lo_hi,
    get_acquire_a_mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380897:4]
  wire  _bundleOut_0_a_valid_T = state == 4'h7; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380901:4]
  wire  _bundleOut_0_a_valid_T_1 = state == 4'h3; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380902:4]
  wire [3:0] get_acquire_size = {{2'd0}, rsize}; // @[Edges.scala 447:17 chipyard.TestHarness.SmallBoomConfig.fir 380827:4 Edges.scala 450:15 chipyard.TestHarness.SmallBoomConfig.fir 380831:4]
  wire  _bundleOut_0_d_ready_T = state == 4'h8; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380921:4]
  wire  _bundleOut_0_d_ready_T_1 = state == 4'h4; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380922:4]
  wire  _T_1 = _io_serial_in_ready_T & io_serial_in_valid; // @[SerialAdapter.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 380929:4]
  wire  _GEN_3 = _T_1 ? 1'h0 : idx; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380930:4 SerialAdapter.scala 140:9 chipyard.TestHarness.SmallBoomConfig.fir 380932:6 SerialAdapter.scala 91:16 chipyard.TestHarness.SmallBoomConfig.fir 380466:4]
  wire [63:0] _GEN_4 = _T_1 ? 64'h0 : addr; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380930:4 SerialAdapter.scala 141:10 chipyard.TestHarness.SmallBoomConfig.fir 380933:6 SerialAdapter.scala 87:17 chipyard.TestHarness.SmallBoomConfig.fir 380462:4]
  wire [63:0] _GEN_5 = _T_1 ? 64'h0 : len; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380930:4 SerialAdapter.scala 142:9 chipyard.TestHarness.SmallBoomConfig.fir 380934:6 SerialAdapter.scala 88:16 chipyard.TestHarness.SmallBoomConfig.fir 380463:4]
  wire [3:0] _GEN_6 = _T_1 ? 4'h1 : state; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380930:4 SerialAdapter.scala 143:11 chipyard.TestHarness.SmallBoomConfig.fir 380935:6 SerialAdapter.scala 97:22 chipyard.TestHarness.SmallBoomConfig.fir 380467:4]
  wire  _T_3 = _io_serial_in_ready_T_1 & io_serial_in_valid; // @[SerialAdapter.scala 146:26 chipyard.TestHarness.SmallBoomConfig.fir 380938:4]
  wire [5:0] _addr_T = {idx,5'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380941:6]
  wire [94:0] _GEN_59 = {{63'd0}, io_serial_in_bits}; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.SmallBoomConfig.fir 380942:6]
  wire [94:0] _addr_T_1 = _GEN_59 << _addr_T; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.SmallBoomConfig.fir 380942:6]
  wire [94:0] _GEN_60 = {{31'd0}, addr}; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 380943:6]
  wire [94:0] _addr_T_2 = _GEN_60 | _addr_T_1; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 380943:6]
  wire  _idx_T_1 = idx + 1'h1; // @[SerialAdapter.scala 148:16 chipyard.TestHarness.SmallBoomConfig.fir 380946:6]
  wire  _GEN_7 = idx ? 1'h0 : _idx_T_1; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.SmallBoomConfig.fir 380949:6 SerialAdapter.scala 150:11 chipyard.TestHarness.SmallBoomConfig.fir 380950:8 SerialAdapter.scala 148:9 chipyard.TestHarness.SmallBoomConfig.fir 380947:6]
  wire [3:0] _GEN_8 = idx ? 4'h2 : _GEN_6; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.SmallBoomConfig.fir 380949:6 SerialAdapter.scala 151:13 chipyard.TestHarness.SmallBoomConfig.fir 380951:8]
  wire [94:0] _GEN_9 = _T_3 ? _addr_T_2 : {{31'd0}, _GEN_4}; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.SmallBoomConfig.fir 380939:4 SerialAdapter.scala 147:10 chipyard.TestHarness.SmallBoomConfig.fir 380944:6]
  wire  _GEN_10 = _T_3 ? _GEN_7 : _GEN_3; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.SmallBoomConfig.fir 380939:4]
  wire [3:0] _GEN_11 = _T_3 ? _GEN_8 : _GEN_6; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.SmallBoomConfig.fir 380939:4]
  wire  _T_6 = _io_serial_in_ready_T_2 & io_serial_in_valid; // @[SerialAdapter.scala 155:25 chipyard.TestHarness.SmallBoomConfig.fir 380955:4]
  wire [94:0] _GEN_62 = {{31'd0}, len}; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.SmallBoomConfig.fir 380960:6]
  wire [94:0] _len_T_2 = _GEN_62 | _addr_T_1; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.SmallBoomConfig.fir 380960:6]
  wire  _T_8 = cmd == 32'h1; // @[SerialAdapter.scala 160:17 chipyard.TestHarness.SmallBoomConfig.fir 380969:8]
  wire  _T_9 = cmd == 32'h0; // @[SerialAdapter.scala 163:24 chipyard.TestHarness.SmallBoomConfig.fir 380975:10]
  wire  _T_12 = ~reset; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.SmallBoomConfig.fir 380982:12]
  wire [3:0] _GEN_12 = _T_9 ? 4'h3 : _GEN_11; // @[SerialAdapter.scala 163:38 chipyard.TestHarness.SmallBoomConfig.fir 380976:10 SerialAdapter.scala 164:15 chipyard.TestHarness.SmallBoomConfig.fir 380977:12]
  wire [1:0] _GEN_13 = _T_8 ? 2'h0 : bodyValid; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.SmallBoomConfig.fir 380970:8 SerialAdapter.scala 161:19 chipyard.TestHarness.SmallBoomConfig.fir 380971:10 SerialAdapter.scala 90:22 chipyard.TestHarness.SmallBoomConfig.fir 380465:4]
  wire [3:0] _GEN_14 = _T_8 ? 4'h6 : _GEN_12; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.SmallBoomConfig.fir 380970:8 SerialAdapter.scala 162:15 chipyard.TestHarness.SmallBoomConfig.fir 380972:10]
  wire  _GEN_15 = idx ? addr[2] : _idx_T_1; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.SmallBoomConfig.fir 380966:6 SerialAdapter.scala 159:11 chipyard.TestHarness.SmallBoomConfig.fir 380968:8 SerialAdapter.scala 157:9 chipyard.TestHarness.SmallBoomConfig.fir 380964:6]
  wire [1:0] _GEN_16 = idx ? _GEN_13 : bodyValid; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.SmallBoomConfig.fir 380966:6 SerialAdapter.scala 90:22 chipyard.TestHarness.SmallBoomConfig.fir 380465:4]
  wire [3:0] _GEN_17 = idx ? _GEN_14 : _GEN_11; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.SmallBoomConfig.fir 380966:6]
  wire [94:0] _GEN_18 = _T_6 ? _len_T_2 : {{31'd0}, _GEN_5}; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.SmallBoomConfig.fir 380956:4 SerialAdapter.scala 156:9 chipyard.TestHarness.SmallBoomConfig.fir 380961:6]
  wire  _GEN_19 = _T_6 ? _GEN_15 : _GEN_10; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.SmallBoomConfig.fir 380956:4]
  wire [1:0] _GEN_20 = _T_6 ? _GEN_16 : bodyValid; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.SmallBoomConfig.fir 380956:4 SerialAdapter.scala 90:22 chipyard.TestHarness.SmallBoomConfig.fir 380465:4]
  wire [3:0] _GEN_21 = _T_6 ? _GEN_17 : _GEN_11; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.SmallBoomConfig.fir 380956:4]
  wire  _T_14 = _bundleOut_0_a_valid_T_1 & auto_out_a_ready; // @[SerialAdapter.scala 171:30 chipyard.TestHarness.SmallBoomConfig.fir 380991:4]
  wire [3:0] _GEN_22 = _T_14 ? 4'h4 : _GEN_21; // @[SerialAdapter.scala 171:46 chipyard.TestHarness.SmallBoomConfig.fir 380992:4 SerialAdapter.scala 172:11 chipyard.TestHarness.SmallBoomConfig.fir 380993:6]
  wire  _T_16 = _bundleOut_0_d_ready_T_1 & auto_out_d_valid; // @[SerialAdapter.scala 175:31 chipyard.TestHarness.SmallBoomConfig.fir 380996:4]
  wire [31:0] _GEN_23 = _T_16 ? auto_out_d_bits_data[31:0] : body_0; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380997:4 SerialAdapter.scala 176:10 chipyard.TestHarness.SmallBoomConfig.fir 381005:6 SerialAdapter.scala 89:17 chipyard.TestHarness.SmallBoomConfig.fir 380464:4]
  wire [31:0] _GEN_24 = _T_16 ? auto_out_d_bits_data[63:32] : body_1; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380997:4 SerialAdapter.scala 176:10 chipyard.TestHarness.SmallBoomConfig.fir 381006:6 SerialAdapter.scala 89:17 chipyard.TestHarness.SmallBoomConfig.fir 380464:4]
  wire  _GEN_25 = _T_16 ? addr[2] : _GEN_19; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380997:4 SerialAdapter.scala 177:9 chipyard.TestHarness.SmallBoomConfig.fir 381008:6]
  wire [94:0] _GEN_26 = _T_16 ? {{63'd0}, nextAddr} : _GEN_9; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380997:4 SerialAdapter.scala 178:10 chipyard.TestHarness.SmallBoomConfig.fir 381009:6]
  wire [3:0] _GEN_27 = _T_16 ? 4'h5 : _GEN_22; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380997:4 SerialAdapter.scala 179:11 chipyard.TestHarness.SmallBoomConfig.fir 381010:6]
  wire  _T_20 = _io_serial_out_valid_T & io_serial_out_ready; // @[SerialAdapter.scala 182:31 chipyard.TestHarness.SmallBoomConfig.fir 381013:4]
  wire [63:0] _len_T_4 = len - 64'h1; // @[SerialAdapter.scala 184:16 chipyard.TestHarness.SmallBoomConfig.fir 381019:6]
  wire  _T_21 = len == 64'h0; // @[SerialAdapter.scala 185:15 chipyard.TestHarness.SmallBoomConfig.fir 381021:6]
  wire [3:0] _GEN_28 = idx ? 4'h3 : _GEN_27; // @[SerialAdapter.scala 186:48 chipyard.TestHarness.SmallBoomConfig.fir 381027:8 SerialAdapter.scala 186:56 chipyard.TestHarness.SmallBoomConfig.fir 381028:10]
  wire [3:0] _GEN_29 = _T_21 ? 4'h0 : _GEN_28; // @[SerialAdapter.scala 185:24 chipyard.TestHarness.SmallBoomConfig.fir 381022:6 SerialAdapter.scala 185:32 chipyard.TestHarness.SmallBoomConfig.fir 381023:8]
  wire  _GEN_30 = _T_20 ? _idx_T_1 : _GEN_25; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.SmallBoomConfig.fir 381014:4 SerialAdapter.scala 183:9 chipyard.TestHarness.SmallBoomConfig.fir 381017:6]
  wire [94:0] _GEN_31 = _T_20 ? {{31'd0}, _len_T_4} : _GEN_18; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.SmallBoomConfig.fir 381014:4 SerialAdapter.scala 184:9 chipyard.TestHarness.SmallBoomConfig.fir 381020:6]
  wire [3:0] _GEN_32 = _T_20 ? _GEN_29 : _GEN_27; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.SmallBoomConfig.fir 381014:4]
  wire  _T_24 = _io_serial_in_ready_T_3 & io_serial_in_valid; // @[SerialAdapter.scala 189:32 chipyard.TestHarness.SmallBoomConfig.fir 381032:4]
  wire [1:0] _bodyValid_T = 2'h1 << idx; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 381035:6]
  wire [1:0] _bodyValid_T_1 = bodyValid | _bodyValid_T; // @[SerialAdapter.scala 191:28 chipyard.TestHarness.SmallBoomConfig.fir 381036:6]
  wire  _T_27 = idx | _T_21; // @[SerialAdapter.scala 192:42 chipyard.TestHarness.SmallBoomConfig.fir 381040:6]
  wire [3:0] _GEN_35 = _T_27 ? 4'h7 : _GEN_32; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.SmallBoomConfig.fir 381041:6 SerialAdapter.scala 193:13 chipyard.TestHarness.SmallBoomConfig.fir 381042:8]
  wire  _GEN_36 = _T_27 ? _GEN_30 : _idx_T_1; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.SmallBoomConfig.fir 381041:6 SerialAdapter.scala 195:11 chipyard.TestHarness.SmallBoomConfig.fir 381047:8]
  wire [94:0] _GEN_37 = _T_27 ? _GEN_31 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.SmallBoomConfig.fir 381041:6 SerialAdapter.scala 196:11 chipyard.TestHarness.SmallBoomConfig.fir 381050:8]
  wire [1:0] _GEN_40 = _T_24 ? _bodyValid_T_1 : _GEN_20; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 381033:4 SerialAdapter.scala 191:15 chipyard.TestHarness.SmallBoomConfig.fir 381037:6]
  wire  _GEN_42 = _T_24 ? _GEN_36 : _GEN_30; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 381033:4]
  wire [94:0] _GEN_43 = _T_24 ? _GEN_37 : _GEN_31; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 381033:4]
  wire  _T_29 = _bundleOut_0_a_valid_T & auto_out_a_ready; // @[SerialAdapter.scala 200:32 chipyard.TestHarness.SmallBoomConfig.fir 381054:4]
  wire  _T_31 = _bundleOut_0_d_ready_T & auto_out_d_valid; // @[SerialAdapter.scala 204:31 chipyard.TestHarness.SmallBoomConfig.fir 381059:4]
  wire [94:0] _GEN_46 = _T_21 ? _GEN_26 : {{63'd0}, nextAddr}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381062:6 SerialAdapter.scala 208:12 chipyard.TestHarness.SmallBoomConfig.fir 381066:8]
  wire [94:0] _GEN_47 = _T_21 ? _GEN_43 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381062:6 SerialAdapter.scala 209:11 chipyard.TestHarness.SmallBoomConfig.fir 381069:8]
  wire  _GEN_48 = _T_21 & _GEN_42; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381062:6 SerialAdapter.scala 210:11 chipyard.TestHarness.SmallBoomConfig.fir 381070:8]
  wire [94:0] _GEN_51 = _T_31 ? _GEN_46 : _GEN_26; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 381060:4]
  wire [94:0] _GEN_52 = _T_31 ? _GEN_47 : _GEN_43; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 381060:4]
  wire  _GEN_67 = _T_6 & idx & ~_T_8 & ~_T_9; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.SmallBoomConfig.fir 380984:14]
  assign auto_out_a_valid = _bundleOut_0_a_valid_T | _bundleOut_0_a_valid_T_1; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380903:4]
  assign auto_out_a_bits_opcode = _bundleOut_0_a_valid_T ? 3'h1 : 3'h4; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380906:4]
  assign auto_out_a_bits_size = _bundleOut_0_a_valid_T ? 4'h3 : get_acquire_size; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380906:4]
  assign auto_out_a_bits_address = _bundleOut_0_a_valid_T ? put_acquire_address : get_acquire_address; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380906:4]
  assign auto_out_a_bits_mask = _bundleOut_0_a_valid_T ? wmask : get_acquire_mask; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380906:4]
  assign auto_out_a_bits_data = _bundleOut_0_a_valid_T ? put_acquire_data : 64'h0; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380906:4]
  assign auto_out_d_ready = _bundleOut_0_d_ready_T | _bundleOut_0_d_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380923:4]
  assign io_serial_in_ready = _io_serial_in_ready_T_5 | _io_serial_in_ready_T_3; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380474:4]
  assign io_serial_out_valid = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.SmallBoomConfig.fir 380476:4]
  assign io_serial_out_bits = idx ? body_1 : body_0; // @[SerialAdapter.scala 101:22 chipyard.TestHarness.SmallBoomConfig.fir 380478:4 SerialAdapter.scala 101:22 chipyard.TestHarness.SmallBoomConfig.fir 380478:4]
  always @(posedge clock) begin
    if (_T_1) begin // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380930:4]
      cmd <= io_serial_in_bits; // @[SerialAdapter.scala 139:9 chipyard.TestHarness.SmallBoomConfig.fir 380931:6]
    end
    addr <= _GEN_51[63:0];
    len <= _GEN_52[63:0];
    if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 381033:4]
      if (~idx) begin // @[SerialAdapter.scala 190:15 chipyard.TestHarness.SmallBoomConfig.fir 381034:6]
        body_0 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.SmallBoomConfig.fir 381034:6]
      end else begin
        body_0 <= _GEN_23;
      end
    end else begin
      body_0 <= _GEN_23;
    end
    if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 381033:4]
      if (idx) begin // @[SerialAdapter.scala 190:15 chipyard.TestHarness.SmallBoomConfig.fir 381034:6]
        body_1 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.SmallBoomConfig.fir 381034:6]
      end else begin
        body_1 <= _GEN_24;
      end
    end else begin
      body_1 <= _GEN_24;
    end
    if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 381060:4]
      if (_T_21) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381062:6]
        bodyValid <= _GEN_40;
      end else begin
        bodyValid <= 2'h0; // @[SerialAdapter.scala 211:17 chipyard.TestHarness.SmallBoomConfig.fir 381071:8]
      end
    end else begin
      bodyValid <= _GEN_40;
    end
    if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 381060:4]
      idx <= _GEN_48;
    end else if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 381033:4]
      if (_T_27) begin // @[SerialAdapter.scala 192:58 chipyard.TestHarness.SmallBoomConfig.fir 381041:6]
        idx <= _GEN_30;
      end else begin
        idx <= _idx_T_1; // @[SerialAdapter.scala 195:11 chipyard.TestHarness.SmallBoomConfig.fir 381047:8]
      end
    end else begin
      idx <= _GEN_30;
    end
    if (reset) begin // @[SerialAdapter.scala 97:22 chipyard.TestHarness.SmallBoomConfig.fir 380467:4]
      state <= 4'h0; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.SmallBoomConfig.fir 380467:4]
    end else if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 381060:4]
      if (_T_21) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381062:6]
        state <= 4'h0; // @[SerialAdapter.scala 206:13 chipyard.TestHarness.SmallBoomConfig.fir 381063:8]
      end else begin
        state <= 4'h6; // @[SerialAdapter.scala 212:13 chipyard.TestHarness.SmallBoomConfig.fir 381072:8]
      end
    end else if (_T_29) begin // @[SerialAdapter.scala 200:48 chipyard.TestHarness.SmallBoomConfig.fir 381055:4]
      state <= 4'h8; // @[SerialAdapter.scala 201:11 chipyard.TestHarness.SmallBoomConfig.fir 381056:6]
    end else if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 381033:4]
      state <= _GEN_35;
    end else begin
      state <= _GEN_32;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & idx & ~_T_8 & ~_T_9 & _T_12) begin
          $fwrite(32'h80000002,
            "Assertion failed: Bad TSI command\n    at SerialAdapter.scala:166 assert(false.B, \"Bad TSI command\")\n"); // @[SerialAdapter.scala 166:15 chipyard.TestHarness.SmallBoomConfig.fir 380984:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_12) begin
          $fatal; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.SmallBoomConfig.fir 380985:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmd = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  len = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  body_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  body_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bodyValid = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  idx = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_53_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 381092:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 381093:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 381094:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input         io_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input         io_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input  [2:0]  io_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 381095:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 383034:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 383341:4]
  wire  _source_ok_T = ~io_in_a_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.SmallBoomConfig.fir 381106:6]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 381111:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 381113:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 381114:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 381114:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 381115:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 381117:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 381118:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 381120:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 381121:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 381122:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 381123:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 381124:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381126:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381127:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381129:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381130:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 381131:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 381132:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 381133:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381134:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381135:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381136:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381137:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381138:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381139:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381140:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381141:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381142:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381143:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381144:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381145:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 381146:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 381147:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 381148:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381149:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381150:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381151:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381152:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381153:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381154:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381155:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381156:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381157:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381158:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381159:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381160:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381161:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381162:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381163:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381164:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381165:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381166:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381167:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381168:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381169:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381170:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381171:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381172:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 381179:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381183:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 381195:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 381198:8]
  wire  _T_20 = _T_17 & _source_ok_T; // @[Parameters.scala 1160:30 chipyard.TestHarness.SmallBoomConfig.fir 381201:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381207:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381208:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381209:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381210:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381212:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381213:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381214:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381215:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381217:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381218:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381219:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381220:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381222:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381223:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h2010000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381224:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381225:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381227:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381228:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381229:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381230:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381232:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381233:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381234:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381235:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381237:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381238:8]
  wire  _T_58 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381239:8]
  wire  _T_65 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48 chipyard.TestHarness.SmallBoomConfig.fir 381246:8]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381248:8]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381249:8]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381251:8]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381252:8]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381253:8]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381254:8]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh10000000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381256:8]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381257:8]
  wire  _T_77 = _T_71 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381258:8]
  wire  _T_78 = _T_65 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381259:8]
  wire  _T_81 = _T_20 & _T_78; // @[Monitor.scala 82:72 chipyard.TestHarness.SmallBoomConfig.fir 381262:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381264:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381265:8]
  wire  _T_147 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381332:8]
  wire  _T_149 = _source_ok_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381338:8]
  wire  _T_150 = ~_T_149; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381339:8]
  wire  _T_153 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381346:8]
  wire  _T_154 = ~_T_153; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381347:8]
  wire  _T_156 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381353:8]
  wire  _T_157 = ~_T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381354:8]
  wire  _T_158 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.SmallBoomConfig.fir 381359:8]
  wire  _T_160 = _T_158 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381361:8]
  wire  _T_161 = ~_T_160; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381362:8]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 381367:8]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 381368:8]
  wire  _T_165 = _T_163 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381370:8]
  wire  _T_166 = ~_T_165; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381371:8]
  wire  _T_167 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.SmallBoomConfig.fir 381376:8]
  wire  _T_169 = _T_167 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381378:8]
  wire  _T_170 = ~_T_169; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381379:8]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 381385:6]
  wire  _T_318 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.SmallBoomConfig.fir 381557:8]
  wire  _T_320 = _T_318 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381559:8]
  wire  _T_321 = ~_T_320; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381560:8]
  wire  _T_331 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 381583:6]
  wire  _T_339 = _T_20 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381592:8]
  wire  _T_340 = ~_T_339; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381593:8]
  wire  _T_350 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381607:8]
  wire  _T_352 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 381609:8]
  wire  _T_395 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381652:8]
  wire  _T_396 = _T_395 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381653:8]
  wire  _T_397 = _T_396 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381654:8]
  wire  _T_398 = _T_397 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381655:8]
  wire  _T_399 = _T_398 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381656:8]
  wire  _T_400 = _T_399 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381657:8]
  wire  _T_401 = _T_400 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381658:8]
  wire  _T_402 = _T_352 & _T_401; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381659:8]
  wire  _T_404 = _T_350 | _T_402; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 381661:8]
  wire  _T_406 = _T_404 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381663:8]
  wire  _T_407 = ~_T_406; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381664:8]
  wire  _T_414 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 381683:8]
  wire  _T_416 = _T_414 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381685:8]
  wire  _T_417 = ~_T_416; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381686:8]
  wire  _T_418 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 381691:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381693:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381694:8]
  wire  _T_426 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 381708:6]
  wire  _T_482 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381765:8]
  wire  _T_483 = _T_482 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381766:8]
  wire  _T_484 = _T_483 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381767:8]
  wire  _T_485 = _T_484 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381768:8]
  wire  _T_486 = _T_485 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381769:8]
  wire  _T_487 = _T_486 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381770:8]
  wire  _T_488 = _T_352 & _T_487; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381771:8]
  wire  _T_497 = _T_350 | _T_488; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 381780:8]
  wire  _T_499 = _T_20 & _T_497; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 381782:8]
  wire  _T_501 = _T_499 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381784:8]
  wire  _T_502 = ~_T_501; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381785:8]
  wire  _T_517 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 381821:6]
  wire [7:0] _T_604 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 381925:8]
  wire [7:0] _T_605 = io_in_a_bits_mask & _T_604; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 381926:8]
  wire  _T_606 = _T_605 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 381927:8]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381929:8]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381930:8]
  wire  _T_610 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 381936:6]
  wire  _T_618 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 381945:8]
  wire  _T_662 = _T_58 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381989:8]
  wire  _T_663 = _T_662 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381990:8]
  wire  _T_664 = _T_663 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381991:8]
  wire  _T_665 = _T_664 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381992:8]
  wire  _T_666 = _T_665 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381993:8]
  wire  _T_667 = _T_666 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381994:8]
  wire  _T_668 = _T_618 & _T_667; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381995:8]
  wire  _T_678 = _T_20 & _T_668; // @[Monitor.scala 131:74 chipyard.TestHarness.SmallBoomConfig.fir 382005:8]
  wire  _T_680 = _T_678 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382007:8]
  wire  _T_681 = ~_T_680; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382008:8]
  wire  _T_688 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.SmallBoomConfig.fir 382027:8]
  wire  _T_690 = _T_688 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382029:8]
  wire  _T_691 = ~_T_690; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382030:8]
  wire  _T_696 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 382044:6]
  wire  _T_774 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.SmallBoomConfig.fir 382135:8]
  wire  _T_776 = _T_774 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382137:8]
  wire  _T_777 = ~_T_776; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382138:8]
  wire  _T_782 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 382152:6]
  wire  _T_851 = _T_352 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 382222:8]
  wire  _T_854 = _T_350 | _T_851; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 382225:8]
  wire  _T_855 = _T_20 & _T_854; // @[Monitor.scala 147:68 chipyard.TestHarness.SmallBoomConfig.fir 382226:8]
  wire  _T_857 = _T_855 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382228:8]
  wire  _T_858 = ~_T_857; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382229:8]
  wire  _T_865 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.SmallBoomConfig.fir 382248:8]
  wire  _T_867 = _T_865 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382250:8]
  wire  _T_868 = ~_T_867; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382251:8]
  wire  _T_877 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 382275:6]
  wire  _T_879 = _T_877 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382277:6]
  wire  _T_880 = ~_T_879; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382278:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.SmallBoomConfig.fir 382283:6]
  wire  _T_881 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 382288:6]
  wire  _T_883 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382291:8]
  wire  _T_884 = ~_T_883; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382292:8]
  wire  _T_885 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 382297:8]
  wire  _T_887 = _T_885 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382299:8]
  wire  _T_888 = ~_T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382300:8]
  wire  _T_889 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.SmallBoomConfig.fir 382305:8]
  wire  _T_891 = _T_889 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382307:8]
  wire  _T_892 = ~_T_891; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382308:8]
  wire  _T_893 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.SmallBoomConfig.fir 382313:8]
  wire  _T_895 = _T_893 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382315:8]
  wire  _T_896 = ~_T_895; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382316:8]
  wire  _T_897 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.SmallBoomConfig.fir 382321:8]
  wire  _T_899 = _T_897 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382323:8]
  wire  _T_900 = ~_T_899; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382324:8]
  wire  _T_901 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 382330:6]
  wire  _T_912 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.SmallBoomConfig.fir 382354:8]
  wire  _T_914 = _T_912 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382356:8]
  wire  _T_915 = ~_T_914; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382357:8]
  wire  _T_916 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.SmallBoomConfig.fir 382362:8]
  wire  _T_918 = _T_916 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382364:8]
  wire  _T_919 = ~_T_918; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382365:8]
  wire  _T_929 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 382388:6]
  wire  _T_949 = _T_897 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.SmallBoomConfig.fir 382429:8]
  wire  _T_951 = _T_949 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382431:8]
  wire  _T_952 = ~_T_951; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382432:8]
  wire  _T_958 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 382447:6]
  wire  _T_975 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 382482:6]
  wire  _T_993 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 382518:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 382584:4]
  wire [8:0] a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 382589:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 382591:4]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382593:4]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 382595:4]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 382596:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 382607:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.SmallBoomConfig.fir 382608:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 382609:4]
  reg  source; // @[Monitor.scala 387:22 chipyard.TestHarness.SmallBoomConfig.fir 382610:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 382611:4]
  wire  _T_1022 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 382612:4]
  wire  _T_1023 = io_in_a_valid & _T_1022; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 382613:4]
  wire  _T_1024 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 382615:6]
  wire  _T_1026 = _T_1024 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382617:6]
  wire  _T_1027 = ~_T_1026; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382618:6]
  wire  _T_1028 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.SmallBoomConfig.fir 382623:6]
  wire  _T_1030 = _T_1028 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382625:6]
  wire  _T_1031 = ~_T_1030; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382626:6]
  wire  _T_1032 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 382631:6]
  wire  _T_1034 = _T_1032 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382633:6]
  wire  _T_1035 = ~_T_1034; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382634:6]
  wire  _T_1036 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.SmallBoomConfig.fir 382639:6]
  wire  _T_1038 = _T_1036 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382641:6]
  wire  _T_1039 = ~_T_1038; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382642:6]
  wire  _T_1040 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 382647:6]
  wire  _T_1042 = _T_1040 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382649:6]
  wire  _T_1043 = ~_T_1042; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382650:6]
  wire  _T_1045 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 382657:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 382665:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 382667:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 382669:4]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 382670:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 382671:4]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382673:4]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 382675:4]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 382676:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 382687:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.SmallBoomConfig.fir 382688:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 382689:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 382690:4]
  reg [2:0] sink; // @[Monitor.scala 539:22 chipyard.TestHarness.SmallBoomConfig.fir 382691:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.SmallBoomConfig.fir 382692:4]
  wire  _T_1046 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 382693:4]
  wire  _T_1047 = io_in_d_valid & _T_1046; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 382694:4]
  wire  _T_1048 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 382696:6]
  wire  _T_1050 = _T_1048 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382698:6]
  wire  _T_1051 = ~_T_1050; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382699:6]
  wire  _T_1052 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.SmallBoomConfig.fir 382704:6]
  wire  _T_1054 = _T_1052 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382706:6]
  wire  _T_1055 = ~_T_1054; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382707:6]
  wire  _T_1056 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 382712:6]
  wire  _T_1058 = _T_1056 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382714:6]
  wire  _T_1059 = ~_T_1058; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382715:6]
  wire  _T_1060 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 382720:6]
  wire  _T_1062 = _T_1060 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382722:6]
  wire  _T_1063 = ~_T_1062; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382723:6]
  wire  _T_1064 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.SmallBoomConfig.fir 382728:6]
  wire  _T_1066 = _T_1064 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382730:6]
  wire  _T_1067 = ~_T_1066; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382731:6]
  wire  _T_1068 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.SmallBoomConfig.fir 382736:6]
  wire  _T_1070 = _T_1068 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382738:6]
  wire  _T_1071 = ~_T_1070; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382739:6]
  wire  _T_1073 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 382746:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 382755:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 382756:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 382757:4]
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382767:4]
  wire [8:0] a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 382769:4]
  wire  a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 382770:4]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382789:4]
  wire [8:0] d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 382791:4]
  wire  d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 382792:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 382813:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 382813:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 382814:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 382818:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 382819:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 382819:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 382820:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.SmallBoomConfig.fir 382824:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 382825:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 382829:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 382830:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 382830:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 382831:4]
  wire  _T_1074 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 382855:4]
  wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 382858:6]
  wire [1:0] _GEN_15 = _T_1074 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 382857:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 382859:6 chipyard.TestHarness.SmallBoomConfig.fir 382806:4]
  wire  _T_1077 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 382862:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 382867:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 382868:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 382870:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 382871:6]
  wire [2:0] _GEN_77 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 382873:6]
  wire [3:0] _a_opcodes_set_T = {{1'd0}, _GEN_77}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 382873:6]
  wire [3:0] a_opcodes_set_interm = _T_1077 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382864:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 382869:6 chipyard.TestHarness.SmallBoomConfig.fir 382852:4]
  wire [18:0] _GEN_78 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 382874:6]
  wire [18:0] _a_opcodes_set_T_1 = _GEN_78 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 382874:6]
  wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 657:77 chipyard.TestHarness.SmallBoomConfig.fir 382876:6]
  wire [4:0] a_sizes_set_interm = _T_1077 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382864:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 382872:6 chipyard.TestHarness.SmallBoomConfig.fir 382854:4]
  wire [19:0] _GEN_79 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 382877:6]
  wire [19:0] _a_sizes_set_T_1 = _GEN_79 << _a_sizes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 382877:6]
  wire  _T_1079 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.SmallBoomConfig.fir 382879:6]
  wire  _T_1081 = ~_T_1079; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 382881:6]
  wire  _T_1083 = _T_1081 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382883:6]
  wire  _T_1084 = ~_T_1083; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382884:6]
  wire [1:0] _GEN_16 = _T_1077 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382864:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 382866:6 chipyard.TestHarness.SmallBoomConfig.fir 382804:4]
  wire [18:0] _GEN_19 = _T_1077 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382864:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 382875:6 chipyard.TestHarness.SmallBoomConfig.fir 382808:4]
  wire [19:0] _GEN_20 = _T_1077 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382864:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 382878:6 chipyard.TestHarness.SmallBoomConfig.fir 382810:4]
  wire  _T_1085 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 382899:4]
  wire  _T_1087 = ~_T_881; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 382901:4]
  wire  _T_1088 = _T_1085 & _T_1087; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 382902:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 382904:6]
  wire [1:0] _GEN_21 = _T_1088 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 382903:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 382905:6 chipyard.TestHarness.SmallBoomConfig.fir 382893:4]
  wire  _T_1090 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 382908:4]
  wire  _T_1093 = _T_1090 & _T_1087; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 382911:4]
  wire [30:0] _GEN_81 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 382920:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_81 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 382920:6]
  wire [30:0] _GEN_82 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.SmallBoomConfig.fir 382927:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_82 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.SmallBoomConfig.fir 382927:6]
  wire [1:0] _GEN_22 = _T_1093 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 382912:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 382914:6 chipyard.TestHarness.SmallBoomConfig.fir 382891:4]
  wire [30:0] _GEN_23 = _T_1093 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 382912:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 382921:6 chipyard.TestHarness.SmallBoomConfig.fir 382895:4]
  wire [30:0] _GEN_24 = _T_1093 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 382912:4 Monitor.scala 678:21 chipyard.TestHarness.SmallBoomConfig.fir 382928:6 chipyard.TestHarness.SmallBoomConfig.fir 382897:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.SmallBoomConfig.fir 382937:6]
  wire  same_cycle_resp = _T_1074 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 382938:6]
  wire  _T_1098 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 382939:6]
  wire  _T_1100 = _T_1098 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 382941:6]
  wire  _T_1102 = _T_1100 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382943:6]
  wire  _T_1103 = ~_T_1102; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382944:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8]
  wire  _T_1104 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382950:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382951:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382951:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382951:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382951:8]
  wire  _T_1105 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382951:8]
  wire  _T_1106 = _T_1104 | _T_1105; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 382952:8]
  wire  _T_1108 = _T_1106 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382954:8]
  wire  _T_1109 = ~_T_1108; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382955:8]
  wire  _T_1110 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 382960:8]
  wire  _T_1112 = _T_1110 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382962:8]
  wire  _T_1113 = ~_T_1112; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382963:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382811:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 382821:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8]
  wire  _T_1115 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382971:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382973:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382973:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382973:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382973:8]
  wire  _T_1117 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382973:8]
  wire  _T_1118 = _T_1115 | _T_1117; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 382974:8]
  wire  _T_1120 = _T_1118 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382976:8]
  wire  _T_1121 = ~_T_1120; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382977:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382822:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 382832:4]
  wire [7:0] _GEN_83 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 382982:8]
  wire  _T_1122 = _GEN_83 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 382982:8]
  wire  _T_1124 = _T_1122 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382984:8]
  wire  _T_1125 = ~_T_1124; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382985:8]
  wire  _T_1127 = _T_1085 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 382993:4]
  wire  _T_1128 = _T_1127 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 382994:4]
  wire  _T_1130 = _T_1128 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 382996:4]
  wire  _T_1132 = _T_1130 & _T_1087; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 382998:4]
  wire  _T_1133 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 383000:6]
  wire  _T_1134 = _T_1133 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 383001:6]
  wire  _T_1136 = _T_1134 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383003:6]
  wire  _T_1137 = ~_T_1136; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383004:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382805:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382892:4]
  wire  _T_1138 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 383010:4]
  wire  _T_1139 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 383011:4]
  wire  _T_1140 = ~_T_1139; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 383012:4]
  wire  _T_1141 = _T_1138 | _T_1140; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 383013:4]
  wire  _T_1143 = _T_1141 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383015:4]
  wire  _T_1144 = ~_T_1143; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383016:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382803:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 383021:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382890:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 383022:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 383023:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382807:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 383025:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382894:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 383026:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 383027:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382809:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 383029:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382896:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.SmallBoomConfig.fir 383030:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 383031:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 383033:4]
  wire  _T_1145 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 383036:4]
  wire  _T_1146 = ~_T_1145; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 383037:4]
  wire  _T_1147 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 383038:4]
  wire  _T_1148 = _T_1146 | _T_1147; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 383039:4]
  wire  _T_1149 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 383040:4]
  wire  _T_1150 = _T_1148 | _T_1149; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 383041:4]
  wire  _T_1152 = _T_1150 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 383043:4]
  wire  _T_1153 = ~_T_1152; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 383044:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 383050:4]
  wire  _T_1156 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 383054:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 383060:4]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383095:4]
  wire [8:0] d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 383097:4]
  wire  d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 383098:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 383131:4]
  wire [15:0] _GEN_87 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 383136:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_87 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 383136:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 383137:4]
  wire  _T_1174 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 383215:4]
  wire  _T_1176 = _T_1174 & _T_881; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 383217:4]
  wire  _T_1178 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 383223:4]
  wire  _T_1180 = _T_1178 & _T_881; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 383225:4]
  wire [30:0] _GEN_69 = _T_1180 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 383226:4 Monitor.scala 786:21 chipyard.TestHarness.SmallBoomConfig.fir 383242:6 chipyard.TestHarness.SmallBoomConfig.fir 383213:4]
  wire  _T_1184 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 383261:6]
  wire  _T_1188 = _T_1184 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383265:6]
  wire  _T_1189 = ~_T_1188; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383266:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 383119:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 383138:4]
  wire  _T_1194 = _GEN_83 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 383284:8]
  wire  _T_1196 = _T_1194 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383286:8]
  wire  _T_1197 = ~_T_1196; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383287:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 383212:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.SmallBoomConfig.fir 383337:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 383338:4]
  wire  _GEN_93 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381267:10]
  wire  _GEN_109 = io_in_a_valid & _T_171; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381457:10]
  wire  _GEN_127 = io_in_a_valid & _T_331; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381595:10]
  wire  _GEN_141 = io_in_a_valid & _T_426; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381787:10]
  wire  _GEN_151 = io_in_a_valid & _T_517; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381900:10]
  wire  _GEN_161 = io_in_a_valid & _T_610; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382010:10]
  wire  _GEN_171 = io_in_a_valid & _T_696; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382118:10]
  wire  _GEN_181 = io_in_a_valid & _T_782; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382231:10]
  wire  _GEN_193 = io_in_d_valid & _T_881; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382294:10]
  wire  _GEN_203 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382336:10]
  wire  _GEN_213 = io_in_d_valid & _T_929; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382394:10]
  wire  _GEN_223 = io_in_d_valid & _T_958; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382453:10]
  wire  _GEN_229 = io_in_d_valid & _T_975; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382488:10]
  wire  _GEN_235 = io_in_d_valid & _T_993; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382524:10]
  wire  _GEN_241 = _T_1088 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382957:10]
  wire  _GEN_246 = _T_1088 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382979:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 383034:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 383341:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382593:4]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382593:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 382603:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 382604:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382592:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382658:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 382659:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382658:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.SmallBoomConfig.fir 382660:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382658:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 382661:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382658:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.SmallBoomConfig.fir 382662:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382658:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 382663:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382673:4]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382673:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 382683:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 382684:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382672:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382747:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 382748:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382747:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.SmallBoomConfig.fir 382749:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382747:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 382750:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382747:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 382751:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382747:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.SmallBoomConfig.fir 382752:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382747:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.SmallBoomConfig.fir 382753:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 382755:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 382755:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 383024:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 382756:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 382756:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 383028:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 382757:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 382757:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 383032:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382767:4]
      a_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382767:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 382777:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 382778:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382592:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382789:4]
      d_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382789:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 382799:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 382800:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382672:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 383033:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 383033:4]
    end else if (_T_1156) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 383055:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 383056:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 383051:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 383060:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 383060:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 383339:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383095:4]
      d_first_counter_2 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383095:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 383105:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 383106:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382672:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381267:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381268:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381334:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381335:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381341:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381342:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381349:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381350:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381356:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381357:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_161) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381364:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_161) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381365:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381373:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381374:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381381:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381382:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381457:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381458:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381524:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381525:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381531:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381532:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381539:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381540:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381546:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381547:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_161) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381554:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_161) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381555:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_321) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381562:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_321) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381563:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381571:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381572:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381579:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381580:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_331 & _T_340) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381595:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_340) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381596:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_407) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381666:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_407) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381667:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381673:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381674:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381680:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381681:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381688:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381689:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381696:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381697:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381704:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381705:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_426 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381787:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381788:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381794:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381795:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381801:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381802:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381809:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381810:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381817:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381818:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_517 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381900:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381901:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381907:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381908:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381914:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381915:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381922:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381923:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381932:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381933:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_610 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382010:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382011:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382017:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382018:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382024:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382025:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_691) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382032:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_691) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382033:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382040:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382041:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_696 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382118:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382119:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382125:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382126:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382132:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382133:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_777) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382140:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_777) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382141:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382148:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382149:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_782 & _T_858) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382231:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_858) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382232:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382238:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382239:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382245:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382246:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_868) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382253:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_868) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382254:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382261:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382262:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382269:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382270:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382280:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382281:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_881 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382294:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382295:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382302:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382303:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382310:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382311:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382318:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382319:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_900) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382326:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_900) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382327:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_901 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382336:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382337:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382351:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382352:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382359:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382360:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382367:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382368:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382375:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382376:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_929 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382394:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382395:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382409:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382410:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382417:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382418:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382425:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382426:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382434:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382435:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_958 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382453:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382454:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382461:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382462:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382469:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382470:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_975 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382488:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382489:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_229 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382496:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382497:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_229 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382505:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382506:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_993 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382524:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382525:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382532:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382533:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382540:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382541:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382620:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382621:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1031) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382628:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1031) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382629:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382636:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382637:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1039) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382644:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1039) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382645:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382652:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382653:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382701:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382702:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382709:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382710:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382717:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382718:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382725:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382726:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382733:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382734:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382741:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382742:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382886:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382887:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382946:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382947:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & same_cycle_resp & _T_1109) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382957:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1109) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382958:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1113) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382965:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1113) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382966:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & ~same_cycle_resp & _T_1121) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382979:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_246 & _T_1121) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382980:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_246 & _T_1125) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382987:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_246 & _T_1125) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382988:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383006:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383007:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1144) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 6 (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383018:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1144) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383019:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1153) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 383046:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1153) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 383047:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383268:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383269:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383289:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383290:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inflight_opcodes = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  inflight_sizes = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerdesser_1_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 383561:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 383562:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 383563:4]
  output        auto_manager_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_manager_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [2:0]  auto_manager_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [2:0]  auto_manager_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [3:0]  auto_manager_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_manager_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [31:0] auto_manager_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [7:0]  auto_manager_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [63:0] auto_manager_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_manager_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_manager_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output        auto_manager_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [2:0]  auto_manager_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [1:0]  auto_manager_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [3:0]  auto_manager_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output        auto_manager_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [2:0]  auto_manager_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output        auto_manager_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [63:0] auto_manager_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output        auto_manager_in_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_client_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output        auto_client_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [2:0]  auto_client_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [2:0]  auto_client_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [2:0]  auto_client_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [3:0]  auto_client_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [28:0] auto_client_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [7:0]  auto_client_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output [63:0] auto_client_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output        auto_client_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output        auto_client_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_client_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [2:0]  auto_client_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [1:0]  auto_client_out_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [2:0]  auto_client_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [3:0]  auto_client_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_client_out_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_client_out_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input  [63:0] auto_client_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  input         auto_client_out_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383564:4]
  output        io_ser_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383565:4]
  input         io_ser_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383565:4]
  input  [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 383565:4]
  input         io_ser_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383565:4]
  output        io_ser_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383565:4]
  output [3:0]  io_ser_out_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 383565:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire [2:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
  wire  outArb_clock; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_reset; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_in_1_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_in_1_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [2:0] outArb_io_in_1_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [2:0] outArb_io_in_1_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [3:0] outArb_io_in_1_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [3:0] outArb_io_in_1_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [63:0] outArb_io_in_1_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_in_1_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [7:0] outArb_io_in_1_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_in_1_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_in_4_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_in_4_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [2:0] outArb_io_in_4_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [2:0] outArb_io_in_4_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [3:0] outArb_io_in_4_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [3:0] outArb_io_in_4_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [31:0] outArb_io_in_4_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [63:0] outArb_io_in_4_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_in_4_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [7:0] outArb_io_in_4_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_in_4_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_out_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_out_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [2:0] outArb_io_out_bits_chanId; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [2:0] outArb_io_out_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [2:0] outArb_io_out_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [3:0] outArb_io_out_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [3:0] outArb_io_out_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [31:0] outArb_io_out_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [63:0] outArb_io_out_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_out_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire [7:0] outArb_io_out_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outArb_io_out_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
  wire  outSer_clock; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire  outSer_reset; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire  outSer_io_in_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire  outSer_io_in_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [2:0] outSer_io_in_bits_chanId; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [2:0] outSer_io_in_bits_opcode; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [2:0] outSer_io_in_bits_param; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [3:0] outSer_io_in_bits_size; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [3:0] outSer_io_in_bits_source; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [31:0] outSer_io_in_bits_address; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [63:0] outSer_io_in_bits_data; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire  outSer_io_in_bits_corrupt; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [7:0] outSer_io_in_bits_union; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire  outSer_io_in_bits_last; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire  outSer_io_out_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire  outSer_io_out_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire [3:0] outSer_io_out_bits; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
  wire  inDes_clock; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire  inDes_reset; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire  inDes_io_in_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire  inDes_io_in_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [3:0] inDes_io_in_bits; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire  inDes_io_out_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire  inDes_io_out_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [2:0] inDes_io_out_bits_chanId; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [2:0] inDes_io_out_bits_opcode; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [2:0] inDes_io_out_bits_param; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [3:0] inDes_io_out_bits_size; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [3:0] inDes_io_out_bits_source; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [31:0] inDes_io_out_bits_address; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [63:0] inDes_io_out_bits_data; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire  inDes_io_out_bits_corrupt; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [7:0] inDes_io_out_bits_union; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
  wire [1:0] _merged_bits_merged_union_T_1 = {auto_client_out_d_bits_sink,auto_client_out_d_bits_denied}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 383664:4]
  wire  merged_1_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383653:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383849:4]
  wire  _merged_bits_last_T_1 = merged_1_ready & auto_client_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 383677:4]
  wire [12:0] _merged_bits_last_beats1_decode_T_1 = 13'h3f << auto_client_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 383679:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_3 = ~_merged_bits_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 383681:4]
  wire [2:0] merged_bits_last_beats1_decode = _merged_bits_last_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 383682:4]
  wire  merged_bits_last_beats1_opdata = auto_client_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 383683:4]
  wire [2:0] merged_bits_last_beats1 = merged_bits_last_beats1_opdata ? merged_bits_last_beats1_decode : 3'h0; // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 383684:4]
  reg [2:0] merged_bits_last_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383685:4]
  wire [2:0] merged_bits_last_counter1_1 = merged_bits_last_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 383687:4]
  wire  merged_bits_last_first_1 = merged_bits_last_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 383688:4]
  wire  _merged_bits_last_last_T_2 = merged_bits_last_counter_1 == 3'h1; // @[Edges.scala 231:25 chipyard.TestHarness.SmallBoomConfig.fir 383689:4]
  wire  _merged_bits_last_last_T_3 = merged_bits_last_beats1 == 3'h0; // @[Edges.scala 231:47 chipyard.TestHarness.SmallBoomConfig.fir 383690:4]
  wire  merged_4_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383796:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383858:4]
  wire  _merged_bits_last_T_4 = merged_4_ready & auto_manager_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 383819:4]
  wire [20:0] _merged_bits_last_beats1_decode_T_13 = 21'h3f << auto_manager_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 383821:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_15 = ~_merged_bits_last_beats1_decode_T_13[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 383823:4]
  wire [2:0] merged_bits_last_beats1_decode_3 = _merged_bits_last_beats1_decode_T_15[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 383824:4]
  wire  merged_bits_last_beats1_opdata_3 = ~auto_manager_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 383826:4]
  wire [2:0] merged_bits_last_beats1_3 = merged_bits_last_beats1_opdata_3 ? merged_bits_last_beats1_decode_3 : 3'h0; // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 383827:4]
  reg [2:0] merged_bits_last_counter_4; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383828:4]
  wire [2:0] merged_bits_last_counter1_4 = merged_bits_last_counter_4 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 383830:4]
  wire  merged_bits_last_first_4 = merged_bits_last_counter_4 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 383831:4]
  wire  _merged_bits_last_last_T_8 = merged_bits_last_counter_4 == 3'h1; // @[Edges.scala 231:25 chipyard.TestHarness.SmallBoomConfig.fir 383832:4]
  wire  _merged_bits_last_last_T_9 = merged_bits_last_beats1_3 == 3'h0; // @[Edges.scala 231:47 chipyard.TestHarness.SmallBoomConfig.fir 383833:4]
  wire  _bundleOut_0_a_valid_T = inDes_io_out_bits_chanId == 3'h0; // @[Serdes.scala 236:37 chipyard.TestHarness.SmallBoomConfig.fir 383871:4]
  wire  _bundleIn_0_d_valid_T = inDes_io_out_bits_chanId == 3'h3; // @[Serdes.scala 239:37 chipyard.TestHarness.SmallBoomConfig.fir 383937:4]
  wire [7:0] _bundleIn_0_d_bits_d_sink_T = {{1'd0}, inDes_io_out_bits_union[7:1]}; // @[Serdes.scala 468:31 chipyard.TestHarness.SmallBoomConfig.fir 383947:4]
  wire  _inDes_io_out_ready_T = 3'h0 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383976:4]
  wire  _inDes_io_out_ready_T_1 = _inDes_io_out_ready_T & auto_client_out_a_ready; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383977:4]
  wire  _inDes_io_out_ready_T_2 = 3'h1 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383978:4]
  wire  _inDes_io_out_ready_T_3 = _inDes_io_out_ready_T_2 ? 1'h0 : _inDes_io_out_ready_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383979:4]
  wire  _inDes_io_out_ready_T_4 = 3'h2 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383980:4]
  wire  _inDes_io_out_ready_T_5 = _inDes_io_out_ready_T_4 ? 1'h0 : _inDes_io_out_ready_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383981:4]
  wire  _inDes_io_out_ready_T_6 = 3'h3 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383982:4]
  wire  _inDes_io_out_ready_T_7 = _inDes_io_out_ready_T_6 ? auto_manager_in_d_ready : _inDes_io_out_ready_T_5; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383983:4]
  wire  _inDes_io_out_ready_T_8 = 3'h4 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383984:4]
  TLMonitor_53_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383575:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  HellaPeekingArbiter_inTestHarness outArb ( // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383606:4]
    .clock(outArb_clock),
    .reset(outArb_reset),
    .io_in_1_ready(outArb_io_in_1_ready),
    .io_in_1_valid(outArb_io_in_1_valid),
    .io_in_1_bits_opcode(outArb_io_in_1_bits_opcode),
    .io_in_1_bits_param(outArb_io_in_1_bits_param),
    .io_in_1_bits_size(outArb_io_in_1_bits_size),
    .io_in_1_bits_source(outArb_io_in_1_bits_source),
    .io_in_1_bits_data(outArb_io_in_1_bits_data),
    .io_in_1_bits_corrupt(outArb_io_in_1_bits_corrupt),
    .io_in_1_bits_union(outArb_io_in_1_bits_union),
    .io_in_1_bits_last(outArb_io_in_1_bits_last),
    .io_in_4_ready(outArb_io_in_4_ready),
    .io_in_4_valid(outArb_io_in_4_valid),
    .io_in_4_bits_opcode(outArb_io_in_4_bits_opcode),
    .io_in_4_bits_param(outArb_io_in_4_bits_param),
    .io_in_4_bits_size(outArb_io_in_4_bits_size),
    .io_in_4_bits_source(outArb_io_in_4_bits_source),
    .io_in_4_bits_address(outArb_io_in_4_bits_address),
    .io_in_4_bits_data(outArb_io_in_4_bits_data),
    .io_in_4_bits_corrupt(outArb_io_in_4_bits_corrupt),
    .io_in_4_bits_union(outArb_io_in_4_bits_union),
    .io_in_4_bits_last(outArb_io_in_4_bits_last),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits_chanId(outArb_io_out_bits_chanId),
    .io_out_bits_opcode(outArb_io_out_bits_opcode),
    .io_out_bits_param(outArb_io_out_bits_param),
    .io_out_bits_size(outArb_io_out_bits_size),
    .io_out_bits_source(outArb_io_out_bits_source),
    .io_out_bits_address(outArb_io_out_bits_address),
    .io_out_bits_data(outArb_io_out_bits_data),
    .io_out_bits_corrupt(outArb_io_out_bits_corrupt),
    .io_out_bits_union(outArb_io_out_bits_union),
    .io_out_bits_last(outArb_io_out_bits_last)
  );
  GenericSerializer_inTestHarness outSer ( // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383609:4]
    .clock(outSer_clock),
    .reset(outSer_reset),
    .io_in_ready(outSer_io_in_ready),
    .io_in_valid(outSer_io_in_valid),
    .io_in_bits_chanId(outSer_io_in_bits_chanId),
    .io_in_bits_opcode(outSer_io_in_bits_opcode),
    .io_in_bits_param(outSer_io_in_bits_param),
    .io_in_bits_size(outSer_io_in_bits_size),
    .io_in_bits_source(outSer_io_in_bits_source),
    .io_in_bits_address(outSer_io_in_bits_address),
    .io_in_bits_data(outSer_io_in_bits_data),
    .io_in_bits_corrupt(outSer_io_in_bits_corrupt),
    .io_in_bits_union(outSer_io_in_bits_union),
    .io_in_bits_last(outSer_io_in_bits_last),
    .io_out_ready(outSer_io_out_ready),
    .io_out_valid(outSer_io_out_valid),
    .io_out_bits(outSer_io_out_bits)
  );
  GenericDeserializer_inTestHarness inDes ( // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383865:4]
    .clock(inDes_clock),
    .reset(inDes_reset),
    .io_in_ready(inDes_io_in_ready),
    .io_in_valid(inDes_io_in_valid),
    .io_in_bits(inDes_io_in_bits),
    .io_out_ready(inDes_io_out_ready),
    .io_out_valid(inDes_io_out_valid),
    .io_out_bits_chanId(inDes_io_out_bits_chanId),
    .io_out_bits_opcode(inDes_io_out_bits_opcode),
    .io_out_bits_param(inDes_io_out_bits_param),
    .io_out_bits_size(inDes_io_out_bits_size),
    .io_out_bits_source(inDes_io_out_bits_source),
    .io_out_bits_address(inDes_io_out_bits_address),
    .io_out_bits_data(inDes_io_out_bits_data),
    .io_out_bits_corrupt(inDes_io_out_bits_corrupt),
    .io_out_bits_union(inDes_io_out_bits_union)
  );
  assign auto_manager_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383796:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383858:4]
  assign auto_manager_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.SmallBoomConfig.fir 383938:4]
  assign auto_manager_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 461:15 chipyard.TestHarness.SmallBoomConfig.fir 383941:4]
  assign auto_manager_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 462:15 chipyard.TestHarness.SmallBoomConfig.fir 383942:4]
  assign auto_manager_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 463:15 chipyard.TestHarness.SmallBoomConfig.fir 383943:4]
  assign auto_manager_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 464:15 chipyard.TestHarness.SmallBoomConfig.fir 383944:4]
  assign auto_manager_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[2:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 468:17 chipyard.TestHarness.SmallBoomConfig.fir 383948:4]
  assign auto_manager_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.SmallBoomConfig.fir 383949:4]
  assign auto_manager_in_d_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 465:15 chipyard.TestHarness.SmallBoomConfig.fir 383945:4]
  assign auto_manager_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 467:17 chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  assign auto_client_out_a_valid = inDes_io_out_valid & _bundleOut_0_a_valid_T; // @[Serdes.scala 631:45 chipyard.TestHarness.SmallBoomConfig.fir 383872:4]
  assign auto_client_out_a_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383874:4 Serdes.scala 375:15 chipyard.TestHarness.SmallBoomConfig.fir 383875:4]
  assign auto_client_out_a_bits_param = inDes_io_out_bits_param; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383874:4 Serdes.scala 376:15 chipyard.TestHarness.SmallBoomConfig.fir 383876:4]
  assign auto_client_out_a_bits_size = inDes_io_out_bits_size[2:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383874:4 Serdes.scala 377:15 chipyard.TestHarness.SmallBoomConfig.fir 383877:4]
  assign auto_client_out_a_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383874:4 Serdes.scala 378:15 chipyard.TestHarness.SmallBoomConfig.fir 383878:4]
  assign auto_client_out_a_bits_address = inDes_io_out_bits_address[28:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383874:4 Serdes.scala 379:15 chipyard.TestHarness.SmallBoomConfig.fir 383879:4]
  assign auto_client_out_a_bits_mask = inDes_io_out_bits_union; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383874:4 Serdes.scala 385:15 chipyard.TestHarness.SmallBoomConfig.fir 383882:4]
  assign auto_client_out_a_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383874:4 Serdes.scala 380:15 chipyard.TestHarness.SmallBoomConfig.fir 383880:4]
  assign auto_client_out_a_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383874:4 Serdes.scala 382:17 chipyard.TestHarness.SmallBoomConfig.fir 383881:4]
  assign auto_client_out_d_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383653:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383849:4]
  assign io_ser_in_ready = inDes_io_in_ready; // @[Serdes.scala 630:17 chipyard.TestHarness.SmallBoomConfig.fir 383870:4]
  assign io_ser_out_valid = outSer_io_out_valid; // @[Serdes.scala 627:16 chipyard.TestHarness.SmallBoomConfig.fir 383863:4]
  assign io_ser_out_bits = outSer_io_out_bits; // @[Serdes.scala 627:16 chipyard.TestHarness.SmallBoomConfig.fir 383862:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 383576:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 383577:4]
  assign monitor_io_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383796:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383858:4]
  assign monitor_io_in_a_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_a_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_a_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_a_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_a_bits_source = auto_manager_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_a_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_a_bits_mask = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_a_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_d_ready = auto_manager_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign monitor_io_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.SmallBoomConfig.fir 383938:4]
  assign monitor_io_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 461:15 chipyard.TestHarness.SmallBoomConfig.fir 383941:4]
  assign monitor_io_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 462:15 chipyard.TestHarness.SmallBoomConfig.fir 383942:4]
  assign monitor_io_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 463:15 chipyard.TestHarness.SmallBoomConfig.fir 383943:4]
  assign monitor_io_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 464:15 chipyard.TestHarness.SmallBoomConfig.fir 383944:4]
  assign monitor_io_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[2:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 468:17 chipyard.TestHarness.SmallBoomConfig.fir 383948:4]
  assign monitor_io_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.SmallBoomConfig.fir 383949:4]
  assign monitor_io_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383940:4 Serdes.scala 467:17 chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  assign outArb_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 383607:4]
  assign outArb_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 383608:4]
  assign outArb_io_in_1_valid = auto_client_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383571:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383598:4]
  assign outArb_io_in_1_bits_opcode = auto_client_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383571:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383598:4]
  assign outArb_io_in_1_bits_param = {{1'd0}, auto_client_out_d_bits_param}; // @[Serdes.scala 312:22 chipyard.TestHarness.SmallBoomConfig.fir 383655:4 Serdes.scala 315:20 chipyard.TestHarness.SmallBoomConfig.fir 383658:4]
  assign outArb_io_in_1_bits_size = {{1'd0}, auto_client_out_d_bits_size}; // @[Serdes.scala 312:22 chipyard.TestHarness.SmallBoomConfig.fir 383655:4 Serdes.scala 316:20 chipyard.TestHarness.SmallBoomConfig.fir 383659:4]
  assign outArb_io_in_1_bits_source = auto_client_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383571:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383598:4]
  assign outArb_io_in_1_bits_data = auto_client_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383571:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383598:4]
  assign outArb_io_in_1_bits_corrupt = auto_client_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383571:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383598:4]
  assign outArb_io_in_1_bits_union = {{6'd0}, _merged_bits_merged_union_T_1}; // @[Serdes.scala 312:22 chipyard.TestHarness.SmallBoomConfig.fir 383655:4 Serdes.scala 322:22 chipyard.TestHarness.SmallBoomConfig.fir 383665:4]
  assign outArb_io_in_1_bits_last = _merged_bits_last_last_T_2 | _merged_bits_last_last_T_3; // @[Edges.scala 231:37 chipyard.TestHarness.SmallBoomConfig.fir 383691:4]
  assign outArb_io_in_4_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign outArb_io_in_4_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign outArb_io_in_4_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign outArb_io_in_4_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign outArb_io_in_4_bits_source = {{3'd0}, auto_manager_in_a_bits_source}; // @[Serdes.scala 255:22 chipyard.TestHarness.SmallBoomConfig.fir 383798:4 Serdes.scala 260:20 chipyard.TestHarness.SmallBoomConfig.fir 383803:4]
  assign outArb_io_in_4_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign outArb_io_in_4_bits_data = auto_manager_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign outArb_io_in_4_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign outArb_io_in_4_bits_union = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383573:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383599:4]
  assign outArb_io_in_4_bits_last = _merged_bits_last_last_T_8 | _merged_bits_last_last_T_9; // @[Edges.scala 231:37 chipyard.TestHarness.SmallBoomConfig.fir 383834:4]
  assign outArb_io_out_ready = outSer_io_in_ready; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383861:4]
  assign outSer_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 383610:4]
  assign outSer_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 383611:4]
  assign outSer_io_in_valid = outArb_io_out_valid; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383860:4]
  assign outSer_io_in_bits_chanId = outArb_io_out_bits_chanId; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_opcode = outArb_io_out_bits_opcode; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_param = outArb_io_out_bits_param; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_size = outArb_io_out_bits_size; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_source = outArb_io_out_bits_source; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_address = outArb_io_out_bits_address; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_data = outArb_io_out_bits_data; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_corrupt = outArb_io_out_bits_corrupt; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_union = outArb_io_out_bits_union; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_in_bits_last = outArb_io_out_bits_last; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383859:4]
  assign outSer_io_out_ready = io_ser_out_ready; // @[Serdes.scala 627:16 chipyard.TestHarness.SmallBoomConfig.fir 383864:4]
  assign inDes_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 383866:4]
  assign inDes_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 383867:4]
  assign inDes_io_in_valid = io_ser_in_valid; // @[Serdes.scala 630:17 chipyard.TestHarness.SmallBoomConfig.fir 383869:4]
  assign inDes_io_in_bits = io_ser_in_bits; // @[Serdes.scala 630:17 chipyard.TestHarness.SmallBoomConfig.fir 383868:4]
  assign inDes_io_out_ready = _inDes_io_out_ready_T_8 ? 1'h0 : _inDes_io_out_ready_T_7; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383985:4]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383685:4]
      merged_bits_last_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383685:4]
    end else if (_merged_bits_last_T_1) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 383695:4]
      if (merged_bits_last_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 383696:6]
        if (merged_bits_last_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 383684:4]
          merged_bits_last_counter_1 <= merged_bits_last_beats1_decode;
        end else begin
          merged_bits_last_counter_1 <= 3'h0;
        end
      end else begin
        merged_bits_last_counter_1 <= merged_bits_last_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383828:4]
      merged_bits_last_counter_4 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383828:4]
    end else if (_merged_bits_last_T_4) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 383838:4]
      if (merged_bits_last_first_4) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 383839:6]
        if (merged_bits_last_beats1_opdata_3) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 383827:4]
          merged_bits_last_counter_4 <= merged_bits_last_beats1_decode_3;
        end else begin
          merged_bits_last_counter_4 <= 3'h0;
        end
      end else begin
        merged_bits_last_counter_4 <= merged_bits_last_counter1_4;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  merged_bits_last_counter_1 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  merged_bits_last_counter_4 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_54_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 384004:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 384005:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 384006:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [7:0]  io_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
  input  [7:0]  io_in_d_bits_source // @[chipyard.TestHarness.SmallBoomConfig.fir 384007:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [159:0] _RAND_10;
  reg [639:0] _RAND_11;
  reg [639:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [159:0] _RAND_16;
  reg [639:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 385498:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 384024:6]
  wire [5:0] _is_aligned_mask_T_1 = 6'h7 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 384030:6]
  wire [2:0] is_aligned_mask = ~_is_aligned_mask_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 384032:6]
  wire [28:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 384033:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 384033:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 384034:6]
  wire [2:0] _mask_sizeOH_T = {{1'd0}, io_in_a_bits_size}; // @[Misc.scala 201:34 chipyard.TestHarness.SmallBoomConfig.fir 384035:6]
  wire [1:0] mask_sizeOH_shiftAmount = _mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 384036:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 384037:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 384039:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 384040:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 384041:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 384042:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 384043:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384045:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384046:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384048:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384049:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 384050:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 384051:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 384052:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384053:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384054:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384055:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384056:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384057:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384058:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384059:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384060:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384061:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384062:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384063:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384064:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 384065:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 384066:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 384067:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384068:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384069:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384070:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384071:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384072:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384073:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384074:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384075:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384076:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384077:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384078:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384079:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384080:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384081:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384082:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384083:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384084:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384085:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384086:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384087:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384088:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384089:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384090:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384091:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 384098:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 384121:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 384137:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 384138:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 384140:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 384141:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384147:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384172:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384173:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384180:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384181:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384187:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384188:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.SmallBoomConfig.fir 384193:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384195:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384196:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 384201:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 384202:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384204:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384205:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.SmallBoomConfig.fir 384210:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384212:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384213:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 384219:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.SmallBoomConfig.fir 384299:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384301:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384302:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 384325:6]
  wire  _T_175 = _T_37 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384359:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384360:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 384379:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384381:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384382:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 384387:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384389:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384390:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 384404:6]
  wire  _T_218 = _source_ok_T_4 & _T_37; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 384430:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384432:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384433:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 384469:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 384525:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 384526:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 384527:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384529:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384530:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 384536:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.SmallBoomConfig.fir 384581:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384583:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384584:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 384598:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.SmallBoomConfig.fir 384643:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384645:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384646:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 384660:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.SmallBoomConfig.fir 384705:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384707:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384708:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 384732:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384734:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384735:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 384746:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 384752:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384755:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384756:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 384761:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384763:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384764:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 384794:6]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 384852:6]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 384911:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 384946:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 384982:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 385048:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385057:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385059:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385060:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 385071:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.SmallBoomConfig.fir 385072:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 385073:4]
  reg [7:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.SmallBoomConfig.fir 385074:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 385075:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 385076:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 385077:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 385079:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385081:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385082:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.SmallBoomConfig.fir 385087:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385089:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385090:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 385095:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385097:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385098:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.SmallBoomConfig.fir 385103:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385105:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385106:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 385111:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385113:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385114:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 385121:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 385129:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385137:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385139:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385140:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 385151:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 385153:4]
  reg [7:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 385154:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 385157:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 385158:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 385160:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385162:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385163:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 385176:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385178:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385179:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 385184:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385186:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385187:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 385210:4]
  reg [159:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 385219:4]
  reg [639:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 385220:4]
  reg [639:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 385221:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385231:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385233:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385234:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385253:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385255:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385256:4]
  wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 385277:4]
  wire [10:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 385277:4]
  wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 385278:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 385282:4]
  wire [639:0] _GEN_73 = {{624'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 385283:4]
  wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 385283:4]
  wire [639:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[639:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 385284:4]
  wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 385289:4]
  wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 385294:4]
  wire [639:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[639:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 385295:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 385319:4]
  wire [255:0] _a_set_wo_ready_T = 256'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 385322:6]
  wire [255:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 385321:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 385323:6 chipyard.TestHarness.SmallBoomConfig.fir 385270:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 385326:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 385331:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 385332:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 385334:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 385335:6]
  wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 385337:6]
  wire [10:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 385337:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385328:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 385333:6 chipyard.TestHarness.SmallBoomConfig.fir 385316:4]
  wire [2050:0] _GEN_79 = {{2047'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 385338:6]
  wire [2050:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 385338:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385328:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 385336:6 chipyard.TestHarness.SmallBoomConfig.fir 385318:4]
  wire [2049:0] _GEN_81 = {{2047'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 385341:6]
  wire [2049:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 385341:6]
  wire [159:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.SmallBoomConfig.fir 385343:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 385345:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385347:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385348:6]
  wire [255:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385328:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 385330:6 chipyard.TestHarness.SmallBoomConfig.fir 385268:4]
  wire [2050:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 2051'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385328:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 385339:6 chipyard.TestHarness.SmallBoomConfig.fir 385272:4]
  wire [2049:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 2050'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385328:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 385342:6 chipyard.TestHarness.SmallBoomConfig.fir 385274:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 385363:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 385365:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 385366:4]
  wire [255:0] _d_clr_wo_ready_T = 256'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 385368:6]
  wire [255:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 385367:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 385369:6 chipyard.TestHarness.SmallBoomConfig.fir 385357:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 385372:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 385375:4]
  wire [2062:0] _GEN_83 = {{2047'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 385384:6]
  wire [2062:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 385384:6]
  wire [255:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 385376:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 385378:6 chipyard.TestHarness.SmallBoomConfig.fir 385355:4]
  wire [2062:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 385376:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 385385:6 chipyard.TestHarness.SmallBoomConfig.fir 385359:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.SmallBoomConfig.fir 385401:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 385402:6]
  wire [159:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 385403:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 385405:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385407:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385408:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385414:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385415:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385415:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385415:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385415:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385415:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 385416:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385418:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385419:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 385424:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385426:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385427:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385275:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 385285:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385435:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385437:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385437:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385437:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385437:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385437:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 385438:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385440:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385441:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385286:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 385296:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 385446:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 385446:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385448:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385449:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 385457:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 385458:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 385460:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 385462:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 385464:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 385465:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385467:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385468:6]
  wire [159:0] a_set_wo_ready = _GEN_15[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385269:4]
  wire [159:0] d_clr_wo_ready = _GEN_21[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385356:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 385474:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 385475:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 385476:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 385477:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385479:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385480:4]
  wire [159:0] a_set = _GEN_16[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385267:4]
  wire [159:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 385485:4]
  wire [159:0] d_clr = _GEN_22[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385354:4]
  wire [159:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 385486:4]
  wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 385487:4]
  wire [639:0] a_opcodes_set = _GEN_19[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385271:4]
  wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 385489:4]
  wire [639:0] d_opcodes_clr = _GEN_23[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385358:4]
  wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 385490:4]
  wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 385491:4]
  wire [639:0] a_sizes_set = _GEN_20[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385273:4]
  wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 385493:4]
  wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 385495:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 385497:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 385500:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 385501:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 385502:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 385503:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 385504:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 385505:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385507:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385508:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 385514:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 385518:4]
  reg [159:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 385522:4]
  reg [639:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 385524:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385559:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385561:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385562:4]
  wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 385595:4]
  wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 385600:4]
  wire [639:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[639:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 385601:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 385679:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 385681:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 385687:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 385689:4]
  wire [255:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 385690:4 Monitor.scala 784:21 chipyard.TestHarness.SmallBoomConfig.fir 385692:6 chipyard.TestHarness.SmallBoomConfig.fir 385671:4]
  wire [2062:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 385690:4 Monitor.scala 785:21 chipyard.TestHarness.SmallBoomConfig.fir 385699:6 chipyard.TestHarness.SmallBoomConfig.fir 385675:4]
  wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 385725:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385729:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385730:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385583:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 385602:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 385748:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385750:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385751:8]
  wire [159:0] d_clr_1 = _GEN_67[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385670:4]
  wire [159:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.SmallBoomConfig.fir 385793:4]
  wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.SmallBoomConfig.fir 385794:4]
  wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385674:4]
  wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.SmallBoomConfig.fir 385797:4]
  wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 385802:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.SmallBoomConfig.fir 385807:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.SmallBoomConfig.fir 385808:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.SmallBoomConfig.fir 385809:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.SmallBoomConfig.fir 385810:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.SmallBoomConfig.fir 385811:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.SmallBoomConfig.fir 385812:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385814:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385815:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.SmallBoomConfig.fir 385821:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384149:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384247:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384344:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384435:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384500:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384564:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384626:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384688:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384758:10]
  wire  _GEN_202 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384800:10]
  wire  _GEN_208 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384858:10]
  wire  _GEN_214 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384917:10]
  wire  _GEN_216 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384952:10]
  wire  _GEN_218 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384988:10]
  wire  _GEN_220 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385421:10]
  wire  _GEN_225 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385443:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 385498:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385057:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385057:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385067:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385068:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385122:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 385123:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385122:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.SmallBoomConfig.fir 385124:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385122:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 385125:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385122:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.SmallBoomConfig.fir 385126:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385122:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 385127:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385137:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385137:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385147:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385148:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 385211:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 385212:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 385211:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 385214:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 385211:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 385215:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 385219:4]
      inflight <= 160'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 385219:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 385488:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 385220:4]
      inflight_opcodes <= 640'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 385220:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 385492:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 385221:4]
      inflight_sizes <= 640'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 385221:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 385496:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385231:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385231:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385241:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385242:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385253:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385253:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385263:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385264:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 385497:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 385497:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 385519:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 385520:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 385515:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 385522:4]
      inflight_1 <= 160'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 385522:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.SmallBoomConfig.fir 385795:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 385524:4]
      inflight_sizes_1 <= 640'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 385524:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 385803:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385559:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385559:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385569:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385570:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.SmallBoomConfig.fir 385828:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.SmallBoomConfig.fir 385829:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.SmallBoomConfig.fir 385822:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384149:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384150:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384168:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384169:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384175:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384176:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384183:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384184:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384190:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384191:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384198:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384199:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384207:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384208:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384215:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384216:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384247:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384248:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384266:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384267:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384273:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384274:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384281:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384282:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384288:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384289:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384296:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384297:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384304:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384305:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384313:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384314:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384321:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384322:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384344:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384345:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384362:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384363:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384369:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384370:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384376:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384377:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384384:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384385:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384392:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384393:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384400:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384401:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384435:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384436:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384442:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384443:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384449:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384450:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384457:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384458:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384465:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384466:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384500:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384501:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384507:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384508:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384514:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384515:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384522:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384523:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384532:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384533:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384564:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384565:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384571:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384572:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384578:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384579:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384586:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384587:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384594:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384595:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384626:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384627:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384633:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384634:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384640:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384641:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384648:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384649:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384656:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384657:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384688:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384689:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384695:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384696:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384702:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384703:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384710:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384711:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384718:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384719:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384726:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384727:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384737:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384738:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384758:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384759:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384766:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384767:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384800:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384801:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384807:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384808:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384815:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384816:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384858:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384859:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384865:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384866:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384873:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384874:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384917:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_214 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384918:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384952:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_216 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384953:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384988:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_218 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384989:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385084:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385085:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385092:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385093:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385100:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385101:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385108:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385109:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385116:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385117:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385165:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385166:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385181:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385182:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385189:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385190:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385350:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385351:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385410:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385411:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385421:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385422:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385429:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385430:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385443:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385444:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385451:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385452:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385470:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385471:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385482:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385483:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385510:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385511:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385732:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385733:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385753:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385754:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385817:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385818:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[7:0];
  _RAND_10 = {5{`RANDOM}};
  inflight = _RAND_10[159:0];
  _RAND_11 = {20{`RANDOM}};
  inflight_opcodes = _RAND_11[639:0];
  _RAND_12 = {20{`RANDOM}};
  inflight_sizes = _RAND_12[639:0];
  _RAND_13 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  watchdog = _RAND_15[31:0];
  _RAND_16 = {5{`RANDOM}};
  inflight_1 = _RAND_16[159:0];
  _RAND_17 = {20{`RANDOM}};
  inflight_sizes_1 = _RAND_17[639:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  watchdog_1 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLRAM_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 385832:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 385833:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 385834:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input  [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input  [7:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  output [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  output [7:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
  output [63:0] auto_in_d_bits_data // @[chipyard.TestHarness.SmallBoomConfig.fir 385835:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [7:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [7:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
  wire [8:0] mem_RW0_addr; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_en; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_clk; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmode; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_wdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_wdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_wdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_wdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_wdata_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_wdata_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_wdata_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_wdata_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_rdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_rdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_rdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_rdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_rdata_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_rdata_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_rdata_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire [7:0] mem_RW0_rdata_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmask_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmask_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmask_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmask_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmask_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmask_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmask_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  wire  mem_RW0_wmask_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
  reg  r_full; // @[SRAM.scala 134:30 chipyard.TestHarness.SmallBoomConfig.fir 385881:4]
  reg [1:0] r_size; // @[SRAM.scala 137:26 chipyard.TestHarness.SmallBoomConfig.fir 385884:4]
  reg [7:0] r_source; // @[SRAM.scala 138:26 chipyard.TestHarness.SmallBoomConfig.fir 385885:4]
  reg  r_read; // @[SRAM.scala 139:26 chipyard.TestHarness.SmallBoomConfig.fir 385886:4]
  reg  REG; // @[SRAM.scala 321:58 chipyard.TestHarness.SmallBoomConfig.fir 386406:4]
  reg [7:0] r_1; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386408:4]
  wire [7:0] r_raw_data_1 = REG ? mem_RW0_rdata_1 : r_1; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386419:4]
  reg [7:0] r_0; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386408:4]
  wire [7:0] r_raw_data_0 = REG ? mem_RW0_rdata_0 : r_0; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386419:4]
  reg [7:0] r_3; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386408:4]
  wire [7:0] r_raw_data_3 = REG ? mem_RW0_rdata_3 : r_3; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386419:4]
  reg [7:0] r_2; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386408:4]
  wire [7:0] r_raw_data_2 = REG ? mem_RW0_rdata_2 : r_2; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386419:4]
  wire [31:0] r_corrected_lo = {r_raw_data_3,r_raw_data_2,r_raw_data_1,r_raw_data_0}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 385949:4]
  reg [7:0] r_5; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386408:4]
  wire [7:0] r_raw_data_5 = REG ? mem_RW0_rdata_5 : r_5; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386419:4]
  reg [7:0] r_4; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386408:4]
  wire [7:0] r_raw_data_4 = REG ? mem_RW0_rdata_4 : r_4; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386419:4]
  reg [7:0] r_7; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386408:4]
  wire [7:0] r_raw_data_7 = REG ? mem_RW0_rdata_7 : r_7; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386419:4]
  reg [7:0] r_6; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386408:4]
  wire [7:0] r_raw_data_6 = REG ? mem_RW0_rdata_6 : r_6; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386419:4]
  wire [31:0] r_corrected_hi = {r_raw_data_7,r_raw_data_6,r_raw_data_5,r_raw_data_4}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 385952:4]
  wire  _bundleIn_0_a_ready_T_2 = ~r_full; // @[SRAM.scala 243:41 chipyard.TestHarness.SmallBoomConfig.fir 386132:4]
  wire  in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.SmallBoomConfig.fir 386133:4]
  wire  a_read = auto_in_a_bits_opcode == 3'h4; // @[SRAM.scala 251:35 chipyard.TestHarness.SmallBoomConfig.fir 386141:4]
  wire  _GEN_22 = auto_in_d_ready ? 1'h0 : r_full; // @[SRAM.scala 273:20 chipyard.TestHarness.SmallBoomConfig.fir 386170:4 SRAM.scala 273:29 chipyard.TestHarness.SmallBoomConfig.fir 386171:6 SRAM.scala 134:30 chipyard.TestHarness.SmallBoomConfig.fir 385881:4]
  wire  _T_18 = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 386173:4]
  wire  _T_19 = ~a_read; // @[SRAM.scala 287:13 chipyard.TestHarness.SmallBoomConfig.fir 386187:6]
  wire  _GEN_24 = _T_18 | _GEN_22; // @[SRAM.scala 274:24 chipyard.TestHarness.SmallBoomConfig.fir 386174:4 SRAM.scala 275:18 chipyard.TestHarness.SmallBoomConfig.fir 386175:6]
  wire  a_lanes_lo_lo_lo = |auto_in_a_bits_mask[0]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386311:4]
  wire  a_lanes_lo_lo_hi = |auto_in_a_bits_mask[1]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386313:4]
  wire  a_lanes_lo_hi_lo = |auto_in_a_bits_mask[2]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386315:4]
  wire  a_lanes_lo_hi_hi = |auto_in_a_bits_mask[3]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386317:4]
  wire  a_lanes_hi_lo_lo = |auto_in_a_bits_mask[4]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386319:4]
  wire  a_lanes_hi_lo_hi = |auto_in_a_bits_mask[5]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386321:4]
  wire  a_lanes_hi_hi_lo = |auto_in_a_bits_mask[6]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386323:4]
  wire  a_lanes_hi_hi_hi = |auto_in_a_bits_mask[7]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386325:4]
  wire [7:0] a_lanes = {a_lanes_hi_hi_hi,a_lanes_hi_hi_lo,a_lanes_hi_lo_hi,a_lanes_hi_lo_lo,a_lanes_lo_hi_hi,
    a_lanes_lo_hi_lo,a_lanes_lo_lo_hi,a_lanes_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 386332:4]
  wire  wen = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.SmallBoomConfig.fir 386340:4]
  wire  _ren_T = ~wen; // @[SRAM.scala 310:15 chipyard.TestHarness.SmallBoomConfig.fir 386343:4]
  wire  ren = _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.SmallBoomConfig.fir 386345:4]
  wire  index_lo_lo_lo = auto_in_a_bits_address[3]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386364:4]
  wire  index_lo_lo_hi = auto_in_a_bits_address[4]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386365:4]
  wire  index_lo_hi_lo = auto_in_a_bits_address[5]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386366:4]
  wire  index_lo_hi_hi = auto_in_a_bits_address[6]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386367:4]
  wire  index_hi_lo_lo = auto_in_a_bits_address[7]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386368:4]
  wire  index_hi_lo_hi = auto_in_a_bits_address[8]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386369:4]
  wire  index_hi_hi_lo = auto_in_a_bits_address[9]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386370:4]
  wire  index_hi_hi_hi_lo = auto_in_a_bits_address[10]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386371:4]
  wire  index_hi_hi_hi_hi = auto_in_a_bits_address[11]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386372:4]
  wire [3:0] index_lo = {index_lo_hi_hi,index_lo_hi_lo,index_lo_lo_hi,index_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 386392:4]
  wire [4:0] index_hi = {index_hi_hi_hi_hi,index_hi_hi_hi_lo,index_hi_hi_lo,index_hi_lo_hi,index_hi_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 386396:4]
  TLMonitor_54_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385842:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source)
  );
  mem_inTestHarness mem ( // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385866:4]
    .RW0_addr(mem_RW0_addr),
    .RW0_en(mem_RW0_en),
    .RW0_clk(mem_RW0_clk),
    .RW0_wmode(mem_RW0_wmode),
    .RW0_wdata_0(mem_RW0_wdata_0),
    .RW0_wdata_1(mem_RW0_wdata_1),
    .RW0_wdata_2(mem_RW0_wdata_2),
    .RW0_wdata_3(mem_RW0_wdata_3),
    .RW0_wdata_4(mem_RW0_wdata_4),
    .RW0_wdata_5(mem_RW0_wdata_5),
    .RW0_wdata_6(mem_RW0_wdata_6),
    .RW0_wdata_7(mem_RW0_wdata_7),
    .RW0_rdata_0(mem_RW0_rdata_0),
    .RW0_rdata_1(mem_RW0_rdata_1),
    .RW0_rdata_2(mem_RW0_rdata_2),
    .RW0_rdata_3(mem_RW0_rdata_3),
    .RW0_rdata_4(mem_RW0_rdata_4),
    .RW0_rdata_5(mem_RW0_rdata_5),
    .RW0_rdata_6(mem_RW0_rdata_6),
    .RW0_rdata_7(mem_RW0_rdata_7),
    .RW0_wmask_0(mem_RW0_wmask_0),
    .RW0_wmask_1(mem_RW0_wmask_1),
    .RW0_wmask_2(mem_RW0_wmask_2),
    .RW0_wmask_3(mem_RW0_wmask_3),
    .RW0_wmask_4(mem_RW0_wmask_4),
    .RW0_wmask_5(mem_RW0_wmask_5),
    .RW0_wmask_6(mem_RW0_wmask_6),
    .RW0_wmask_7(mem_RW0_wmask_7)
  );
  assign auto_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.SmallBoomConfig.fir 386133:4]
  assign auto_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.SmallBoomConfig.fir 386112:4]
  assign auto_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 SRAM.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 386060:4]
  assign auto_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.SmallBoomConfig.fir 386062:4]
  assign auto_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.SmallBoomConfig.fir 386064:4]
  assign auto_in_d_bits_data = {r_corrected_hi,r_corrected_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 385960:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 385843:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 385844:4]
  assign monitor_io_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.SmallBoomConfig.fir 386133:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385865:4]
  assign monitor_io_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.SmallBoomConfig.fir 386112:4]
  assign monitor_io_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385840:4 SRAM.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 386060:4]
  assign monitor_io_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.SmallBoomConfig.fir 386062:4]
  assign monitor_io_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.SmallBoomConfig.fir 386064:4]
  assign mem_RW0_wdata_0 = auto_in_a_bits_data[7:0]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386192:4]
  assign mem_RW0_wdata_1 = auto_in_a_bits_data[15:8]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386193:4]
  assign mem_RW0_wdata_2 = auto_in_a_bits_data[23:16]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386194:4]
  assign mem_RW0_wdata_3 = auto_in_a_bits_data[31:24]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386195:4]
  assign mem_RW0_wdata_4 = auto_in_a_bits_data[39:32]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386196:4]
  assign mem_RW0_wdata_5 = auto_in_a_bits_data[47:40]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386197:4]
  assign mem_RW0_wdata_6 = auto_in_a_bits_data[55:48]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386198:4]
  assign mem_RW0_wdata_7 = auto_in_a_bits_data[63:56]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386199:4]
  assign mem_RW0_wmask_0 = a_lanes[0]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386429:6]
  assign mem_RW0_wmask_1 = a_lanes[1]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386430:6]
  assign mem_RW0_wmask_2 = a_lanes[2]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386431:6]
  assign mem_RW0_wmask_3 = a_lanes[3]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386432:6]
  assign mem_RW0_wmask_4 = a_lanes[4]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386433:6]
  assign mem_RW0_wmask_5 = a_lanes[5]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386434:6]
  assign mem_RW0_wmask_6 = a_lanes[6]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386435:6]
  assign mem_RW0_wmask_7 = a_lanes[7]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386436:6]
  assign mem_RW0_wmode = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.SmallBoomConfig.fir 386340:4]
  assign mem_RW0_clk = clock;
  assign mem_RW0_en = ren | wen;
  assign mem_RW0_addr = {index_hi,index_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 386397:4]
  always @(posedge clock) begin
    if (reset) begin // @[SRAM.scala 134:30 chipyard.TestHarness.SmallBoomConfig.fir 385881:4]
      r_full <= 1'h0; // @[SRAM.scala 134:30 chipyard.TestHarness.SmallBoomConfig.fir 385881:4]
    end else begin
      r_full <= _GEN_24;
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.SmallBoomConfig.fir 386174:4]
      r_size <= auto_in_a_bits_size; // @[SRAM.scala 279:18 chipyard.TestHarness.SmallBoomConfig.fir 386179:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.SmallBoomConfig.fir 386174:4]
      r_source <= auto_in_a_bits_source; // @[SRAM.scala 280:18 chipyard.TestHarness.SmallBoomConfig.fir 386180:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.SmallBoomConfig.fir 386174:4]
      r_read <= a_read; // @[SRAM.scala 281:18 chipyard.TestHarness.SmallBoomConfig.fir 386181:6]
    end
    REG <= _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.SmallBoomConfig.fir 386345:4]
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386409:4]
      r_1 <= mem_RW0_rdata_1; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386411:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386409:4]
      r_0 <= mem_RW0_rdata_0; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386410:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386409:4]
      r_3 <= mem_RW0_rdata_3; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386413:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386409:4]
      r_2 <= mem_RW0_rdata_2; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386412:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386409:4]
      r_5 <= mem_RW0_rdata_5; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386415:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386409:4]
      r_4 <= mem_RW0_rdata_4; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386414:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386409:4]
      r_7 <= mem_RW0_rdata_7; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386417:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386409:4]
      r_6 <= mem_RW0_rdata_6; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386416:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_size = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  r_source = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  r_read = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  r_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  r_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  r_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  r_5 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  r_4 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  r_7 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  r_6 = _RAND_12[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar_10_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 386473:2]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [3:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [3:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [2:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [3:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [2:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [3:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 386476:4]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386481:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386485:4]
  assign auto_in_d_valid = auto_out_d_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.SmallBoomConfig.fir 386897:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386481:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386485:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386481:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386485:4]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386481:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386485:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Xbar.scala 228:69 chipyard.TestHarness.SmallBoomConfig.fir 386596:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Xbar.scala 323:53 chipyard.TestHarness.SmallBoomConfig.fir 386658:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386481:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386485:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386481:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386485:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386481:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386485:4]
  assign auto_out_a_valid = auto_in_a_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.SmallBoomConfig.fir 386922:4]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386483:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386486:4]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386483:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386486:4]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386483:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386486:4]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55 chipyard.TestHarness.SmallBoomConfig.fir 386550:4]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386483:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386486:4]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386483:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386486:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386483:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386486:4]
  assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386483:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386486:4]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386483:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386486:4]
endmodule
module TLMonitor_55_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 386999:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 387000:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 387001:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [7:0]  io_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input  [7:0]  io_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 387002:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [159:0] _RAND_13;
  reg [639:0] _RAND_14;
  reg [639:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [159:0] _RAND_19;
  reg [639:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 388493:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 388800:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 387019:6]
  wire [5:0] _is_aligned_mask_T_1 = 6'h7 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 387025:6]
  wire [2:0] is_aligned_mask = ~_is_aligned_mask_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 387027:6]
  wire [28:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 387028:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 387028:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 387029:6]
  wire [2:0] _mask_sizeOH_T = {{1'd0}, io_in_a_bits_size}; // @[Misc.scala 201:34 chipyard.TestHarness.SmallBoomConfig.fir 387030:6]
  wire [1:0] mask_sizeOH_shiftAmount = _mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 387031:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 387032:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 387034:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 387035:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 387036:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 387037:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 387038:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387040:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387041:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387043:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387044:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 387045:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 387046:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 387047:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387048:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387049:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387050:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387051:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387052:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387053:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387054:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387055:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387056:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387057:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387058:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387059:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 387060:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 387061:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 387062:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387063:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387064:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387065:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387066:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387067:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387068:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387069:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387070:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387071:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387072:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387073:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387074:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387075:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387076:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387077:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387078:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387079:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387080:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387081:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387082:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387083:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387084:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387085:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387086:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 387093:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 387116:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 387132:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 387133:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 387135:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 387136:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387142:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387167:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387168:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387175:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387176:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387182:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387183:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.SmallBoomConfig.fir 387188:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387190:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387191:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 387196:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 387197:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387199:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387200:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.SmallBoomConfig.fir 387205:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387207:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387208:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 387214:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.SmallBoomConfig.fir 387294:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387296:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387297:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 387320:6]
  wire  _T_175 = _T_37 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387354:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387355:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 387374:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387376:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387377:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 387382:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387384:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387385:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 387399:6]
  wire  _T_218 = _source_ok_T_4 & _T_37; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 387425:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387427:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387428:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 387464:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 387520:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 387521:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 387522:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387524:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387525:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 387531:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.SmallBoomConfig.fir 387576:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387578:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387579:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 387593:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.SmallBoomConfig.fir 387638:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387640:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387641:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 387655:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.SmallBoomConfig.fir 387700:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387702:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387703:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 387727:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387729:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387730:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 387741:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 387747:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387750:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387751:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 387756:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387758:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387759:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.SmallBoomConfig.fir 387764:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387766:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387767:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.SmallBoomConfig.fir 387772:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387774:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387775:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.SmallBoomConfig.fir 387780:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387782:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387783:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 387789:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.SmallBoomConfig.fir 387813:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387815:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387816:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.SmallBoomConfig.fir 387821:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387823:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387824:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 387847:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.SmallBoomConfig.fir 387888:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387890:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387891:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 387906:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 387941:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 387977:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 388043:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388052:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388054:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388055:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 388066:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.SmallBoomConfig.fir 388067:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 388068:4]
  reg [7:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.SmallBoomConfig.fir 388069:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 388070:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 388071:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 388072:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 388074:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388076:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388077:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.SmallBoomConfig.fir 388082:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388084:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388085:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 388090:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388092:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388093:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.SmallBoomConfig.fir 388098:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388100:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388101:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 388106:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388108:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388109:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 388116:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 388124:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388132:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388134:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388135:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 388146:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.SmallBoomConfig.fir 388147:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 388148:4]
  reg [7:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 388149:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.SmallBoomConfig.fir 388150:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.SmallBoomConfig.fir 388151:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 388152:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 388153:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 388155:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388157:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388158:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.SmallBoomConfig.fir 388163:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388165:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388166:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 388171:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388173:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388174:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 388179:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388181:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388182:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.SmallBoomConfig.fir 388187:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388189:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388190:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.SmallBoomConfig.fir 388195:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388197:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388198:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 388205:4]
  reg [159:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 388214:4]
  reg [639:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 388215:4]
  reg [639:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 388216:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388226:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388228:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388229:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388248:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388250:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388251:4]
  wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 388272:4]
  wire [10:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 388272:4]
  wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 388273:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 388277:4]
  wire [639:0] _GEN_73 = {{624'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 388278:4]
  wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 388278:4]
  wire [639:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[639:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 388279:4]
  wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 388284:4]
  wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 388289:4]
  wire [639:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[639:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 388290:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 388314:4]
  wire [255:0] _a_set_wo_ready_T = 256'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 388317:6]
  wire [255:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 388316:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 388318:6 chipyard.TestHarness.SmallBoomConfig.fir 388265:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 388321:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 388326:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 388327:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 388329:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 388330:6]
  wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 388332:6]
  wire [10:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 388332:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388323:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 388328:6 chipyard.TestHarness.SmallBoomConfig.fir 388311:4]
  wire [2050:0] _GEN_79 = {{2047'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 388333:6]
  wire [2050:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 388333:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388323:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 388331:6 chipyard.TestHarness.SmallBoomConfig.fir 388313:4]
  wire [2049:0] _GEN_81 = {{2047'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 388336:6]
  wire [2049:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 388336:6]
  wire [159:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.SmallBoomConfig.fir 388338:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 388340:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388342:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388343:6]
  wire [255:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388323:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 388325:6 chipyard.TestHarness.SmallBoomConfig.fir 388263:4]
  wire [2050:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 2051'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388323:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 388334:6 chipyard.TestHarness.SmallBoomConfig.fir 388267:4]
  wire [2049:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 2050'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388323:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 388337:6 chipyard.TestHarness.SmallBoomConfig.fir 388269:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 388358:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 388360:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 388361:4]
  wire [255:0] _d_clr_wo_ready_T = 256'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 388363:6]
  wire [255:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 388362:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 388364:6 chipyard.TestHarness.SmallBoomConfig.fir 388352:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 388367:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 388370:4]
  wire [2062:0] _GEN_83 = {{2047'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 388379:6]
  wire [2062:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 388379:6]
  wire [255:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 388371:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 388373:6 chipyard.TestHarness.SmallBoomConfig.fir 388350:4]
  wire [2062:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 388371:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 388380:6 chipyard.TestHarness.SmallBoomConfig.fir 388354:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.SmallBoomConfig.fir 388396:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 388397:6]
  wire [159:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 388398:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 388400:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388402:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388403:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388409:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388410:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388410:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388410:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388410:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388410:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 388411:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388413:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388414:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 388419:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388421:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388422:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388270:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 388280:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388430:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388432:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388432:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388432:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388432:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388432:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 388433:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388435:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388436:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388281:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 388291:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 388441:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 388441:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388443:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388444:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 388452:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 388453:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 388455:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 388457:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 388459:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 388460:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388462:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388463:6]
  wire [159:0] a_set_wo_ready = _GEN_15[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388264:4]
  wire [159:0] d_clr_wo_ready = _GEN_21[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388351:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 388469:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 388470:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 388471:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 388472:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388474:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388475:4]
  wire [159:0] a_set = _GEN_16[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388262:4]
  wire [159:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 388480:4]
  wire [159:0] d_clr = _GEN_22[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388349:4]
  wire [159:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 388481:4]
  wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 388482:4]
  wire [639:0] a_opcodes_set = _GEN_19[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388266:4]
  wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 388484:4]
  wire [639:0] d_opcodes_clr = _GEN_23[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388353:4]
  wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 388485:4]
  wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 388486:4]
  wire [639:0] a_sizes_set = _GEN_20[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388268:4]
  wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 388488:4]
  wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 388490:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 388492:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 388495:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 388496:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 388497:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 388498:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 388499:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 388500:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388502:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388503:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 388509:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 388513:4]
  reg [159:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 388517:4]
  reg [639:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 388519:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388554:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388556:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388557:4]
  wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 388590:4]
  wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 388595:4]
  wire [639:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[639:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 388596:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 388674:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 388676:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 388682:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 388684:4]
  wire [255:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 388685:4 Monitor.scala 784:21 chipyard.TestHarness.SmallBoomConfig.fir 388687:6 chipyard.TestHarness.SmallBoomConfig.fir 388666:4]
  wire [2062:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 388685:4 Monitor.scala 785:21 chipyard.TestHarness.SmallBoomConfig.fir 388694:6 chipyard.TestHarness.SmallBoomConfig.fir 388670:4]
  wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 388720:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388724:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388725:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388578:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 388597:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 388743:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388745:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388746:8]
  wire [159:0] d_clr_1 = _GEN_67[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388665:4]
  wire [159:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.SmallBoomConfig.fir 388788:4]
  wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.SmallBoomConfig.fir 388789:4]
  wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388669:4]
  wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.SmallBoomConfig.fir 388792:4]
  wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 388797:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 388799:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.SmallBoomConfig.fir 388802:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.SmallBoomConfig.fir 388803:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.SmallBoomConfig.fir 388804:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.SmallBoomConfig.fir 388805:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.SmallBoomConfig.fir 388806:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.SmallBoomConfig.fir 388807:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388809:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388810:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.SmallBoomConfig.fir 388816:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387144:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387242:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387339:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387430:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387495:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387559:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387621:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387683:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387753:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387795:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387853:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387912:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387947:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387983:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388416:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388438:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 388493:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 388800:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388052:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388052:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388062:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388063:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388117:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 388118:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388117:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.SmallBoomConfig.fir 388119:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388117:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 388120:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388117:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.SmallBoomConfig.fir 388121:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388117:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 388122:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388132:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388132:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388142:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388143:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388206:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 388207:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388206:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.SmallBoomConfig.fir 388208:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388206:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 388209:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388206:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 388210:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388206:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.SmallBoomConfig.fir 388211:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388206:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.SmallBoomConfig.fir 388212:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 388214:4]
      inflight <= 160'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 388214:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 388483:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 388215:4]
      inflight_opcodes <= 640'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 388215:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 388487:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 388216:4]
      inflight_sizes <= 640'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 388216:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 388491:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388226:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388226:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388236:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388237:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388248:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388248:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388258:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388259:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 388492:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 388492:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 388514:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 388515:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 388510:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 388517:4]
      inflight_1 <= 160'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 388517:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.SmallBoomConfig.fir 388790:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 388519:4]
      inflight_sizes_1 <= 640'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 388519:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 388798:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388554:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388554:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388564:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388565:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 388799:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 388799:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.SmallBoomConfig.fir 388823:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.SmallBoomConfig.fir 388824:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.SmallBoomConfig.fir 388817:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387144:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387145:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387163:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387164:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387170:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387171:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387178:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387179:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387185:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387186:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387193:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387194:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387202:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387203:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387210:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387211:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387242:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387243:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387261:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387262:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387268:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387269:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387276:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387277:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387283:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387284:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387291:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387292:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387299:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387300:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387308:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387309:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387316:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387317:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387339:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387340:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387357:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387358:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387364:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387365:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387371:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387372:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387379:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387380:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387387:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387388:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387395:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387396:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387430:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387431:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387437:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387438:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387444:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387445:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387452:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387453:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387460:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387461:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387495:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387496:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387502:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387503:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387509:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387510:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387517:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387518:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387527:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387528:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387559:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387560:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387566:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387567:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387573:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387574:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387581:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387582:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387589:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387590:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387621:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387622:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387628:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387629:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387635:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387636:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387643:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387644:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387651:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387652:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387683:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387684:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387690:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387691:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387697:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387698:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387705:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387706:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387713:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387714:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387721:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387722:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387732:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387733:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387753:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387754:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387761:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387762:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387769:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387770:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387777:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387778:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387785:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387786:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387795:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387796:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387802:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387803:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387810:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387811:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387818:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387819:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387826:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387827:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387834:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387835:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387843:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387844:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387853:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387854:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387860:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387861:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387868:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387869:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387876:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387877:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387884:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387885:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387893:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387894:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387902:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387903:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387912:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387913:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387920:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387921:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387928:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387929:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387937:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387938:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387947:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387948:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387955:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387956:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387964:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387965:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387973:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387974:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387983:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387984:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387991:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387992:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387999:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388000:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388008:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388009:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388079:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388080:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388087:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388088:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388095:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388096:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388103:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388104:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388111:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388112:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388160:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388161:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388168:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388169:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388176:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388177:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388184:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388185:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388192:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388193:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388200:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388201:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388345:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388346:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388405:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388406:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388416:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388417:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388424:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388425:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388438:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388439:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388446:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388447:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388465:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388466:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388477:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388478:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388505:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388506:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388727:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388728:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388748:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388749:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388812:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388813:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {5{`RANDOM}};
  inflight = _RAND_13[159:0];
  _RAND_14 = {20{`RANDOM}};
  inflight_opcodes = _RAND_14[639:0];
  _RAND_15 = {20{`RANDOM}};
  inflight_sizes = _RAND_15[639:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {5{`RANDOM}};
  inflight_1 = _RAND_19[159:0];
  _RAND_20 = {20{`RANDOM}};
  inflight_sizes_1 = _RAND_20[639:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_44_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 388827:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 388828:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 388829:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input  [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input  [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input  [7:0]  io_enq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input  [28:0] io_enq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output [7:0]  io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output [28:0] io_deq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 388830:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  reg [7:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [7:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [7:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  reg [28:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [28:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [28:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388833:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388834:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 388835:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 388836:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 388837:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 388838:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 388839:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 388840:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 388843:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 388858:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 388864:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 388867:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 388873:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 388871:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388883:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388882:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388881:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388880:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388879:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388878:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388877:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388876:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388832:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388833:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388833:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 388846:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 388859:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388834:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388834:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 388861:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 388865:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 388835:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 388835:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 388868:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 388869:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[28:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_20_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 388955:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 388956:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 388957:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [7:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [7:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [7:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [7:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  input  [63:0] auto_out_d_bits_data // @[chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [7:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire [7:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [1:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [28:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire  bundleOut_0_a_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [1:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [28:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [7:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [7:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire  bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
  TLMonitor_55_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388965:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_44_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388992:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_5_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 389006:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 389004:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 389005:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 389018:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 388966:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 388967:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 389004:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 389019:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 388993:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 388994:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388990:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 389007:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 389008:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388990:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388990:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388990:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388990:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388988:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388990:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388963:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388991:4]
endmodule
module TLMonitor_56_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 389055:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 389056:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 389057:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [2:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [3:0]  io_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [2:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input  [3:0]  io_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 389058:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 390549:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 390856:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 4'h9; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 389075:6]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 389081:6]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 389083:6]
  wire [28:0] _GEN_71 = {{23'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 389084:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 389084:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 389085:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 389087:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 389088:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 389090:6]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 389091:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 389092:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 389093:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 389094:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389096:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389097:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389099:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389100:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 389101:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 389102:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 389103:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389104:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389105:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389106:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389107:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389108:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389109:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389110:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389111:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389112:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389113:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389114:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389115:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 389116:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 389117:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 389118:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389119:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389120:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389121:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389122:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389123:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389124:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389125:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389126:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389127:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389128:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389129:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389130:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389131:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389132:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389133:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389134:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389135:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389136:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389137:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389138:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389139:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389140:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389141:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389142:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 389149:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 389172:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 389188:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 389189:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 389191:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 389192:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389198:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389223:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389224:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389231:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389232:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389238:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389239:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.SmallBoomConfig.fir 389244:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389246:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389247:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 389252:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 389253:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389255:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389256:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.SmallBoomConfig.fir 389261:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389263:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389264:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 389270:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.SmallBoomConfig.fir 389350:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389352:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389353:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 389376:6]
  wire  _T_164 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 389399:8]
  wire  _T_172 = _T_164 & _T_37; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 389407:8]
  wire  _T_175 = _T_172 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389410:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389411:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 389430:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389432:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389433:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 389438:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389440:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389441:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 389455:6]
  wire  _T_218 = _source_ok_T_4 & _T_172; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 389481:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389483:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389484:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 389520:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 389576:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 389577:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 389578:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389580:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389581:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 389587:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.SmallBoomConfig.fir 389632:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389634:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389635:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 389649:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.SmallBoomConfig.fir 389694:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389696:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389697:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 389711:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.SmallBoomConfig.fir 389756:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389758:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389759:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 389783:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389785:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389786:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 4'h9; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 389797:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 389803:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389806:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389807:8]
  wire  _T_405 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 389812:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389814:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389815:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.SmallBoomConfig.fir 389820:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389822:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389823:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.SmallBoomConfig.fir 389828:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389830:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389831:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.SmallBoomConfig.fir 389836:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389838:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389839:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 389845:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.SmallBoomConfig.fir 389869:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389871:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389872:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.SmallBoomConfig.fir 389877:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389879:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389880:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 389903:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.SmallBoomConfig.fir 389944:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389946:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389947:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 389962:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 389997:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 390033:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390099:4]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 390104:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 390106:4]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390108:4]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390110:4]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390111:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 390122:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.SmallBoomConfig.fir 390123:4]
  reg [2:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 390124:4]
  reg [3:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.SmallBoomConfig.fir 390125:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 390126:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 390127:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 390128:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 390130:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390132:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390133:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.SmallBoomConfig.fir 390138:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390140:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390141:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 390146:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390148:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390149:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.SmallBoomConfig.fir 390154:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390156:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390157:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 390162:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390164:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390165:6]
  wire  _T_565 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 390172:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390180:4]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 390182:4]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 390184:4]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 390185:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 390186:4]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390188:4]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390190:4]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390191:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 390202:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.SmallBoomConfig.fir 390203:4]
  reg [2:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 390204:4]
  reg [3:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 390205:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.SmallBoomConfig.fir 390206:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.SmallBoomConfig.fir 390207:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 390208:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 390209:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 390211:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390213:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390214:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.SmallBoomConfig.fir 390219:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390221:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390222:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 390227:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390229:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390230:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 390235:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390237:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390238:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.SmallBoomConfig.fir 390243:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390245:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390246:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.SmallBoomConfig.fir 390251:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390253:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390254:6]
  wire  _T_593 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 390261:4]
  reg [9:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 390270:4]
  reg [39:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 390271:4]
  reg [39:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 390272:4]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390282:4]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390284:4]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390285:4]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390304:4]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390306:4]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390307:4]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 390328:4]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 390328:4]
  wire [39:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 390329:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 390333:4]
  wire [39:0] _GEN_73 = {{24'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 390334:4]
  wire [39:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 390334:4]
  wire [39:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[39:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 390335:4]
  wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 390340:4]
  wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 390345:4]
  wire [39:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[39:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 390346:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 390370:4]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 390373:6]
  wire [15:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 390372:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 390374:6 chipyard.TestHarness.SmallBoomConfig.fir 390321:4]
  wire  _T_597 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 390377:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 390382:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 390383:6]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 390385:6]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 390386:6]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 390388:6]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 390388:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390379:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 390384:6 chipyard.TestHarness.SmallBoomConfig.fir 390367:4]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 390389:6]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 390389:6]
  wire [3:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390379:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 390387:6 chipyard.TestHarness.SmallBoomConfig.fir 390369:4]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 390392:6]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 390392:6]
  wire [9:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.SmallBoomConfig.fir 390394:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 390396:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390398:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390399:6]
  wire [15:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390379:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 390381:6 chipyard.TestHarness.SmallBoomConfig.fir 390319:4]
  wire [130:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390379:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 390390:6 chipyard.TestHarness.SmallBoomConfig.fir 390323:4]
  wire [130:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390379:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 390393:6 chipyard.TestHarness.SmallBoomConfig.fir 390325:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 390414:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 390416:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 390417:4]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 390419:6]
  wire [15:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 390418:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 390420:6 chipyard.TestHarness.SmallBoomConfig.fir 390408:4]
  wire  _T_610 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 390423:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 390426:4]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 390435:6]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 390435:6]
  wire [15:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 390427:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 390429:6 chipyard.TestHarness.SmallBoomConfig.fir 390406:4]
  wire [142:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 390427:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 390436:6 chipyard.TestHarness.SmallBoomConfig.fir 390410:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.SmallBoomConfig.fir 390452:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 390453:6]
  wire [9:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 390454:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 390456:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390458:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390459:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390465:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390466:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390466:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390466:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390466:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390466:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 390467:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390469:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390470:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 390475:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390477:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390478:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390326:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 390336:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390486:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390488:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390488:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390488:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390488:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390488:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 390489:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390491:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390492:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390337:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 390347:4]
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 390497:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 390497:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390499:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390500:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 390508:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 390509:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 390511:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 390513:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 390515:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 390516:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390518:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390519:6]
  wire [9:0] a_set_wo_ready = _GEN_15[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390320:4]
  wire [9:0] d_clr_wo_ready = _GEN_21[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390407:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 390525:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 390526:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 390527:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 390528:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390530:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390531:4]
  wire [9:0] a_set = _GEN_16[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390318:4]
  wire [9:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 390536:4]
  wire [9:0] d_clr = _GEN_22[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390405:4]
  wire [9:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 390537:4]
  wire [9:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 390538:4]
  wire [39:0] a_opcodes_set = _GEN_19[39:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390322:4]
  wire [39:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 390540:4]
  wire [39:0] d_opcodes_clr = _GEN_23[39:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390409:4]
  wire [39:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 390541:4]
  wire [39:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 390542:4]
  wire [39:0] a_sizes_set = _GEN_20[39:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390324:4]
  wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 390544:4]
  wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 390546:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 390548:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 390551:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 390552:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 390553:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 390554:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 390555:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 390556:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390558:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390559:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 390565:4]
  wire  _T_676 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 390569:4]
  reg [9:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 390573:4]
  reg [39:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 390575:4]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390610:4]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390612:4]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390613:4]
  wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 390646:4]
  wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 390651:4]
  wire [39:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[39:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 390652:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 390730:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 390732:4]
  wire  _T_698 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 390738:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 390740:4]
  wire [15:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 390741:4 Monitor.scala 784:21 chipyard.TestHarness.SmallBoomConfig.fir 390743:6 chipyard.TestHarness.SmallBoomConfig.fir 390722:4]
  wire [142:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 390741:4 Monitor.scala 785:21 chipyard.TestHarness.SmallBoomConfig.fir 390750:6 chipyard.TestHarness.SmallBoomConfig.fir 390726:4]
  wire [9:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 390776:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390780:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390781:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390634:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 390653:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 390799:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390801:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390802:8]
  wire [9:0] d_clr_1 = _GEN_67[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390721:4]
  wire [9:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.SmallBoomConfig.fir 390844:4]
  wire [9:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.SmallBoomConfig.fir 390845:4]
  wire [39:0] d_opcodes_clr_1 = _GEN_68[39:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390725:4]
  wire [39:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.SmallBoomConfig.fir 390848:4]
  wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 390853:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 390855:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.SmallBoomConfig.fir 390858:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.SmallBoomConfig.fir 390859:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.SmallBoomConfig.fir 390860:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.SmallBoomConfig.fir 390861:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.SmallBoomConfig.fir 390862:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.SmallBoomConfig.fir 390863:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390865:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390866:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.SmallBoomConfig.fir 390872:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389200:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389298:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389395:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389486:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389551:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389615:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389677:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389739:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389809:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389851:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389909:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389968:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390003:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390039:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390472:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390494:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 390549:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 390856:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390108:4]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390108:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390118:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390119:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390107:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390173:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 390174:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390173:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.SmallBoomConfig.fir 390175:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390173:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 390176:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390173:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.SmallBoomConfig.fir 390177:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390173:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 390178:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390188:4]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390188:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390198:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390199:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390187:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390262:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 390263:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390262:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.SmallBoomConfig.fir 390264:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390262:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 390265:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390262:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 390266:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390262:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.SmallBoomConfig.fir 390267:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390262:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.SmallBoomConfig.fir 390268:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 390270:4]
      inflight <= 10'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 390270:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 390539:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 390271:4]
      inflight_opcodes <= 40'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 390271:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 390543:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 390272:4]
      inflight_sizes <= 40'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 390272:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 390547:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390282:4]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390282:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390292:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390293:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390107:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390304:4]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390304:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390314:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390315:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390187:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 390548:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 390548:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 390570:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 390571:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 390566:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 390573:4]
      inflight_1 <= 10'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 390573:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.SmallBoomConfig.fir 390846:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 390575:4]
      inflight_sizes_1 <= 40'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 390575:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 390854:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390610:4]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390610:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390620:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390621:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390187:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 390855:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 390855:4]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47 chipyard.TestHarness.SmallBoomConfig.fir 390879:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.SmallBoomConfig.fir 390880:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.SmallBoomConfig.fir 390873:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389200:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389201:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389219:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389220:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389226:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389227:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389234:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389235:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389241:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389242:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389249:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389250:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389258:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389259:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389266:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389267:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389298:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389299:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389317:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389318:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389324:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389325:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389332:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389333:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389339:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389340:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389347:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389348:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389355:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389356:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389364:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389365:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389372:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389373:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389395:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389396:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389413:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389414:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389420:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389421:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389427:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389428:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389435:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389436:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389443:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389444:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389451:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389452:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389486:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389487:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389493:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389494:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389500:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389501:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389508:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389509:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389516:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389517:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389551:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389552:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389558:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389559:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389565:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389566:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389573:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389574:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389583:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389584:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389615:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389616:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389622:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389623:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389629:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389630:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389637:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389638:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389645:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389646:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389677:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389678:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389684:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389685:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389691:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389692:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389699:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389700:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389707:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389708:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389739:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389740:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389746:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389747:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389753:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389754:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389761:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389762:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389769:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389770:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389777:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389778:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389788:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389789:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389809:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389810:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389817:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389818:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389825:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389826:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389833:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389834:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389841:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389842:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389851:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389852:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389858:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389859:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389866:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389867:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389874:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389875:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389882:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389883:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389890:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389891:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389899:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389900:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389909:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389910:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389916:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389917:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389924:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389925:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389932:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389933:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389940:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389941:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389949:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389950:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389958:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389959:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389968:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389969:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389976:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389977:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389984:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389985:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389993:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389994:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390003:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390004:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390011:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390012:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390020:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390021:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390029:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390030:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390039:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390040:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390047:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390048:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390055:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390056:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390064:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390065:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390135:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390136:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390143:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390144:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390151:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390152:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390159:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390160:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390167:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390168:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390216:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390217:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390224:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390225:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390232:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390233:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390240:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390241:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390248:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390249:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390256:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390257:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390401:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390402:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390461:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390462:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390472:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390473:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390480:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390481:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390494:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390495:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390502:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390503:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390521:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390522:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390533:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390534:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390561:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390562:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390783:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390784:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390804:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390805:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390868:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390869:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[9:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_opcodes = _RAND_14[39:0];
  _RAND_15 = {2{`RANDOM}};
  inflight_sizes = _RAND_15[39:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_1 = _RAND_19[9:0];
  _RAND_20 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_20[39:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_7_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 390883:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 390884:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 390885:4]
  input         io_repeat, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output        io_full, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input  [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input  [2:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input  [3:0]  io_enq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input  [28:0] io_enq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output [2:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output [3:0]  io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output [28:0] io_deq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 390886:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21 chipyard.TestHarness.SmallBoomConfig.fir 390888:4]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390889:4]
  reg [2:0] saved_param; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390889:4]
  reg [2:0] saved_size; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390889:4]
  reg [3:0] saved_source; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390889:4]
  reg [28:0] saved_address; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390889:4]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390889:4]
  reg  saved_corrupt; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390889:4]
  wire  _io_enq_ready_T = ~full; // @[Repeater.scala 24:35 chipyard.TestHarness.SmallBoomConfig.fir 390892:4]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390905:4]
  wire  _T_1 = _T & io_repeat; // @[Repeater.scala 28:23 chipyard.TestHarness.SmallBoomConfig.fir 390906:4]
  wire  _GEN_0 = _T_1 | full; // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390907:4 Repeater.scala 28:45 chipyard.TestHarness.SmallBoomConfig.fir 390908:6 Repeater.scala 19:21 chipyard.TestHarness.SmallBoomConfig.fir 390888:4]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390918:4]
  wire  _T_3 = ~io_repeat; // @[Repeater.scala 29:26 chipyard.TestHarness.SmallBoomConfig.fir 390919:4]
  wire  _T_4 = _T_2 & _T_3; // @[Repeater.scala 29:23 chipyard.TestHarness.SmallBoomConfig.fir 390920:4]
  assign io_full = full; // @[Repeater.scala 26:11 chipyard.TestHarness.SmallBoomConfig.fir 390904:4]
  assign io_enq_ready = io_deq_ready & _io_enq_ready_T; // @[Repeater.scala 24:32 chipyard.TestHarness.SmallBoomConfig.fir 390893:4]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32 chipyard.TestHarness.SmallBoomConfig.fir 390890:4]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390895:4]
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390895:4]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390895:4]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390895:4]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390895:4]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390895:4]
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390895:4]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21 chipyard.TestHarness.SmallBoomConfig.fir 390888:4]
      full <= 1'h0; // @[Repeater.scala 19:21 chipyard.TestHarness.SmallBoomConfig.fir 390888:4]
    end else if (_T_4) begin // @[Repeater.scala 29:38 chipyard.TestHarness.SmallBoomConfig.fir 390921:4]
      full <= 1'h0; // @[Repeater.scala 29:45 chipyard.TestHarness.SmallBoomConfig.fir 390922:6]
    end else begin
      full <= _GEN_0;
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390907:4]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390916:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390907:4]
      saved_param <= io_enq_bits_param; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390915:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390907:4]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390914:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390907:4]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390913:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390907:4]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390912:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390907:4]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390911:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390907:4]
      saved_corrupt <= io_enq_bits_corrupt; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390909:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  saved_mask = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  saved_corrupt = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_7_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 390925:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 390926:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 390927:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [3:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [3:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [7:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [7:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 390928:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire  repeater_clock; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_reset; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [2:0] repeater_io_enq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [3:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [28:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_io_enq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [2:0] repeater_io_deq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [3:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [28:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  wire  repeater_io_deq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29 chipyard.TestHarness.SmallBoomConfig.fir 390962:4]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24 chipyard.TestHarness.SmallBoomConfig.fir 390963:4]
  reg  dToggle; // @[Fragmenter.scala 191:30 chipyard.TestHarness.SmallBoomConfig.fir 390964:4]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41 chipyard.TestHarness.SmallBoomConfig.fir 390965:4]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29 chipyard.TestHarness.SmallBoomConfig.fir 390966:4]
  wire  dLast = dFragnum == 3'h0; // @[Fragmenter.scala 194:30 chipyard.TestHarness.SmallBoomConfig.fir 390967:4]
  wire [3:0] dsizeOH = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 390969:4]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 390972:4]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 390974:4]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 390975:4]
  wire  ack_decrement = dHasData | dsizeOH[3]; // @[Fragmenter.scala 204:32 chipyard.TestHarness.SmallBoomConfig.fir 390992:4]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47 chipyard.TestHarness.SmallBoomConfig.fir 390993:4]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69 chipyard.TestHarness.SmallBoomConfig.fir 390994:4]
  wire [5:0] dFirst_size_lo = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69 chipyard.TestHarness.SmallBoomConfig.fir 390994:4]
  wire [6:0] _dFirst_size_T_1 = {dFirst_size_lo, 1'h0}; // @[package.scala 232:35 chipyard.TestHarness.SmallBoomConfig.fir 390995:4]
  wire [6:0] _dFirst_size_T_2 = _dFirst_size_T_1 | 7'h1; // @[package.scala 232:40 chipyard.TestHarness.SmallBoomConfig.fir 390996:4]
  wire [6:0] _dFirst_size_T_3 = {1'h0,dFirst_size_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 390997:4]
  wire [6:0] _dFirst_size_T_4 = ~_dFirst_size_T_3; // @[package.scala 232:53 chipyard.TestHarness.SmallBoomConfig.fir 390998:4]
  wire [6:0] _dFirst_size_T_5 = _dFirst_size_T_2 & _dFirst_size_T_4; // @[package.scala 232:51 chipyard.TestHarness.SmallBoomConfig.fir 390999:4]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_5[6:4]; // @[OneHot.scala 30:18 chipyard.TestHarness.SmallBoomConfig.fir 391000:4]
  wire [3:0] dFirst_size_lo_1 = _dFirst_size_T_5[3:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.SmallBoomConfig.fir 391001:4]
  wire  dFirst_size_hi_1 = |dFirst_size_hi; // @[OneHot.scala 32:14 chipyard.TestHarness.SmallBoomConfig.fir 391002:4]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28 chipyard.TestHarness.SmallBoomConfig.fir 391003:4]
  wire [3:0] _dFirst_size_T_6 = _GEN_8 | dFirst_size_lo_1; // @[OneHot.scala 32:28 chipyard.TestHarness.SmallBoomConfig.fir 391003:4]
  wire [1:0] dFirst_size_hi_2 = _dFirst_size_T_6[3:2]; // @[OneHot.scala 30:18 chipyard.TestHarness.SmallBoomConfig.fir 391004:4]
  wire [1:0] dFirst_size_lo_2 = _dFirst_size_T_6[1:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.SmallBoomConfig.fir 391005:4]
  wire  dFirst_size_hi_3 = |dFirst_size_hi_2; // @[OneHot.scala 32:14 chipyard.TestHarness.SmallBoomConfig.fir 391006:4]
  wire [1:0] _dFirst_size_T_7 = dFirst_size_hi_2 | dFirst_size_lo_2; // @[OneHot.scala 32:28 chipyard.TestHarness.SmallBoomConfig.fir 391007:4]
  wire  dFirst_size_lo_3 = _dFirst_size_T_7[1]; // @[CircuitMath.scala 30:8 chipyard.TestHarness.SmallBoomConfig.fir 391008:4]
  wire [2:0] dFirst_size = {dFirst_size_hi_1,dFirst_size_hi_3,dFirst_size_lo_3}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 391010:4]
  wire  _drop_T = ~dHasData; // @[Fragmenter.scala 222:20 chipyard.TestHarness.SmallBoomConfig.fir 391023:4]
  wire  _drop_T_2 = ~dLast; // @[Fragmenter.scala 222:33 chipyard.TestHarness.SmallBoomConfig.fir 391025:4]
  wire  drop = _drop_T & _drop_T_2; // @[Fragmenter.scala 222:30 chipyard.TestHarness.SmallBoomConfig.fir 391026:4]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.SmallBoomConfig.fir 391027:4]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 391011:4]
  wire [2:0] _GEN_9 = {{2'd0}, ack_decrement}; // @[Fragmenter.scala 209:55 chipyard.TestHarness.SmallBoomConfig.fir 391013:6]
  wire [2:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55 chipyard.TestHarness.SmallBoomConfig.fir 391014:6]
  wire  _bundleIn_0_d_valid_T = ~drop; // @[Fragmenter.scala 224:39 chipyard.TestHarness.SmallBoomConfig.fir 391029:4]
  wire  _aFrag_T = repeater_io_deq_bits_size > 3'h3; // @[Fragmenter.scala 285:31 chipyard.TestHarness.SmallBoomConfig.fir 391062:4]
  wire [2:0] aFrag = _aFrag_T ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24 chipyard.TestHarness.SmallBoomConfig.fir 391063:4]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 391065:4]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 391067:4]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 391069:4]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 391071:4]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 391073:4]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29 chipyard.TestHarness.SmallBoomConfig.fir 391075:4]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29 chipyard.TestHarness.SmallBoomConfig.fir 391076:4]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79 chipyard.TestHarness.SmallBoomConfig.fir 391079:4]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30 chipyard.TestHarness.SmallBoomConfig.fir 391080:4]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28 chipyard.TestHarness.SmallBoomConfig.fir 391081:4]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26 chipyard.TestHarness.SmallBoomConfig.fir 391084:4]
  reg  aToggle_r; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 391091:4]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 391092:4 Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 391093:6 Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 391091:4]
  wire  bundleOut_0_a_bits_source_hi_lo = ~_GEN_5; // @[Fragmenter.scala 297:23 chipyard.TestHarness.SmallBoomConfig.fir 391096:4]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391105:4]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 391097:4]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31 chipyard.TestHarness.SmallBoomConfig.fir 391101:4]
  wire  _repeater_io_repeat_T_1 = new_gennum != 3'h0; // @[Fragmenter.scala 302:53 chipyard.TestHarness.SmallBoomConfig.fir 391102:4]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65 chipyard.TestHarness.SmallBoomConfig.fir 391106:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90 chipyard.TestHarness.SmallBoomConfig.fir 391107:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88 chipyard.TestHarness.SmallBoomConfig.fir 391108:4]
  wire [5:0] _GEN_10 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100 chipyard.TestHarness.SmallBoomConfig.fir 391109:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100 chipyard.TestHarness.SmallBoomConfig.fir 391109:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111 chipyard.TestHarness.SmallBoomConfig.fir 391110:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51 chipyard.TestHarness.SmallBoomConfig.fir 391111:4]
  wire [28:0] _GEN_11 = {{23'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49 chipyard.TestHarness.SmallBoomConfig.fir 391112:4]
  wire [4:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,bundleOut_0_a_bits_source_hi_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 391114:4]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17 chipyard.TestHarness.SmallBoomConfig.fir 391118:4]
  wire  _T_11 = _T_9 | _repeater_io_repeat_T; // @[Fragmenter.scala 309:35 chipyard.TestHarness.SmallBoomConfig.fir 391120:4]
  wire  _T_13 = _T_11 | reset; // @[Fragmenter.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 391122:4]
  wire  _T_14 = ~_T_13; // @[Fragmenter.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 391123:4]
  wire  _T_16 = repeater_io_deq_bits_mask == 8'hff; // @[Fragmenter.scala 312:53 chipyard.TestHarness.SmallBoomConfig.fir 391130:4]
  wire  _T_17 = _T_9 | _T_16; // @[Fragmenter.scala 312:35 chipyard.TestHarness.SmallBoomConfig.fir 391131:4]
  wire  _T_19 = _T_17 | reset; // @[Fragmenter.scala 312:16 chipyard.TestHarness.SmallBoomConfig.fir 391133:4]
  wire  _T_20 = ~_T_19; // @[Fragmenter.scala 312:16 chipyard.TestHarness.SmallBoomConfig.fir 391134:4]
  TLMonitor_56_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Repeater_7_inTestHarness repeater ( // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_param(repeater_io_enq_bits_param),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_param(repeater_io_deq_bits_param),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 Fragmenter.scala 263:25 chipyard.TestHarness.SmallBoomConfig.fir 391041:4]
  assign auto_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.SmallBoomConfig.fir 391030:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.SmallBoomConfig.fir 391035:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source[7:4]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.SmallBoomConfig.fir 391033:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391105:4]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391105:4]
  assign auto_out_a_bits_param = repeater_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391105:4]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 Fragmenter.scala 306:25 chipyard.TestHarness.SmallBoomConfig.fir 391117:4]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 391115:4]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49 chipyard.TestHarness.SmallBoomConfig.fir 391112:4]
  assign auto_out_a_bits_mask = repeater_io_full ? 8'hff : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31 chipyard.TestHarness.SmallBoomConfig.fir 391139:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391105:4]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.SmallBoomConfig.fir 391027:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 390936:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 390937:4]
  assign monitor_io_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 Fragmenter.scala 263:25 chipyard.TestHarness.SmallBoomConfig.fir 391041:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign monitor_io_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.SmallBoomConfig.fir 391030:4]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign monitor_io_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.SmallBoomConfig.fir 391035:4]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:4]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.SmallBoomConfig.fir 391033:4]
  assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  assign repeater_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 391039:4]
  assign repeater_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 391040:4]
  assign repeater_io_repeat = _repeater_io_repeat_T & _repeater_io_repeat_T_1; // @[Fragmenter.scala 302:41 chipyard.TestHarness.SmallBoomConfig.fir 391103:4]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign repeater_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390933:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390961:4]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390958:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390960:4]
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29 chipyard.TestHarness.SmallBoomConfig.fir 390962:4]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29 chipyard.TestHarness.SmallBoomConfig.fir 390962:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.SmallBoomConfig.fir 391012:4]
      if (dFirst) begin // @[Fragmenter.scala 209:24 chipyard.TestHarness.SmallBoomConfig.fir 391015:6]
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.SmallBoomConfig.fir 391012:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.SmallBoomConfig.fir 391017:6]
        dOrig <= dFirst_size; // @[Fragmenter.scala 211:19 chipyard.TestHarness.SmallBoomConfig.fir 391018:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30 chipyard.TestHarness.SmallBoomConfig.fir 390964:4]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30 chipyard.TestHarness.SmallBoomConfig.fir 390964:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.SmallBoomConfig.fir 391012:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.SmallBoomConfig.fir 391017:6]
        dToggle <= auto_out_d_bits_source[3]; // @[Fragmenter.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 391020:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29 chipyard.TestHarness.SmallBoomConfig.fir 391075:4]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29 chipyard.TestHarness.SmallBoomConfig.fir 391075:4]
    end else if (_T_8) begin // @[Fragmenter.scala 300:29 chipyard.TestHarness.SmallBoomConfig.fir 391098:4]
      gennum <= new_gennum; // @[Fragmenter.scala 300:38 chipyard.TestHarness.SmallBoomConfig.fir 391099:6]
    end
    if (aFirst) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 391092:4]
      aToggle_r <= dToggle; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 391093:6]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 391125:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_14) begin
          $fatal; // @[Fragmenter.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 391126:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16 chipyard.TestHarness.SmallBoomConfig.fir 391136:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_20) begin
          $fatal; // @[Fragmenter.scala 312:16 chipyard.TestHarness.SmallBoomConfig.fir 391137:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_57_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 391177:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 391178:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 391179:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input  [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input  [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input  [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input         io_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input  [2:0]  io_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 391180:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 393119:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 393426:4]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 391196:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 391198:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 391199:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 391199:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 391200:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 391202:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 391203:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 391205:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 391206:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 391207:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 391208:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 391209:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391211:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391212:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391214:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391215:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 391216:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 391217:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 391218:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391219:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391220:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391221:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391222:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391223:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391224:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391225:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391226:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391227:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391228:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391229:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391230:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 391231:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 391232:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 391233:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391234:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391235:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391236:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391237:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391238:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391239:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391240:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391241:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391242:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391243:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391244:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391245:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391246:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391247:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391248:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391249:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391250:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391251:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391252:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391253:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391254:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391255:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391256:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391257:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 391264:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391268:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 391280:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 391283:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391292:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391293:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391294:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391295:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391297:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391298:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391299:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391300:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391302:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391303:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391304:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391305:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391307:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391308:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h2010000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391309:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391310:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391312:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391313:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391314:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391315:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391317:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391318:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391319:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391320:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391322:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391323:8]
  wire  _T_58 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391324:8]
  wire  _T_65 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48 chipyard.TestHarness.SmallBoomConfig.fir 391331:8]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391333:8]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391334:8]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391336:8]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391337:8]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391338:8]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391339:8]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh10000000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391341:8]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391342:8]
  wire  _T_77 = _T_71 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391343:8]
  wire  _T_78 = _T_65 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 391344:8]
  wire  _T_81 = _T_17 & _T_78; // @[Monitor.scala 82:72 chipyard.TestHarness.SmallBoomConfig.fir 391347:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391349:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391350:8]
  wire  _T_147 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391417:8]
  wire  _T_153 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391431:8]
  wire  _T_154 = ~_T_153; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391432:8]
  wire  _T_156 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391438:8]
  wire  _T_157 = ~_T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391439:8]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 391452:8]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 391453:8]
  wire  _T_165 = _T_163 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391455:8]
  wire  _T_166 = ~_T_165; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391456:8]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 391470:6]
  wire  _T_331 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 391668:6]
  wire  _T_339 = _T_17 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391677:8]
  wire  _T_340 = ~_T_339; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391678:8]
  wire  _T_350 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 391692:8]
  wire  _T_352 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 391694:8]
  wire  _T_395 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391737:8]
  wire  _T_396 = _T_395 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391738:8]
  wire  _T_397 = _T_396 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391739:8]
  wire  _T_398 = _T_397 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391740:8]
  wire  _T_399 = _T_398 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391741:8]
  wire  _T_400 = _T_399 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391742:8]
  wire  _T_401 = _T_400 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391743:8]
  wire  _T_402 = _T_352 & _T_401; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 391744:8]
  wire  _T_404 = _T_350 | _T_402; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 391746:8]
  wire  _T_406 = _T_404 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391748:8]
  wire  _T_407 = ~_T_406; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391749:8]
  wire  _T_418 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 391776:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391778:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391779:8]
  wire  _T_426 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 391793:6]
  wire  _T_482 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391850:8]
  wire  _T_483 = _T_482 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391851:8]
  wire  _T_484 = _T_483 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391852:8]
  wire  _T_485 = _T_484 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391853:8]
  wire  _T_486 = _T_485 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391854:8]
  wire  _T_487 = _T_486 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391855:8]
  wire  _T_488 = _T_352 & _T_487; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 391856:8]
  wire  _T_497 = _T_350 | _T_488; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 391865:8]
  wire  _T_499 = _T_17 & _T_497; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 391867:8]
  wire  _T_501 = _T_499 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391869:8]
  wire  _T_502 = ~_T_501; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391870:8]
  wire  _T_517 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 391906:6]
  wire [7:0] _T_604 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 392010:8]
  wire [7:0] _T_605 = io_in_a_bits_mask & _T_604; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 392011:8]
  wire  _T_606 = _T_605 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 392012:8]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392014:8]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392015:8]
  wire  _T_610 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 392021:6]
  wire  _T_618 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 392030:8]
  wire  _T_662 = _T_58 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392074:8]
  wire  _T_663 = _T_662 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392075:8]
  wire  _T_664 = _T_663 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392076:8]
  wire  _T_665 = _T_664 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392077:8]
  wire  _T_666 = _T_665 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392078:8]
  wire  _T_667 = _T_666 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392079:8]
  wire  _T_668 = _T_618 & _T_667; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 392080:8]
  wire  _T_678 = _T_17 & _T_668; // @[Monitor.scala 131:74 chipyard.TestHarness.SmallBoomConfig.fir 392090:8]
  wire  _T_680 = _T_678 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392092:8]
  wire  _T_681 = ~_T_680; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392093:8]
  wire  _T_696 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 392129:6]
  wire  _T_782 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 392237:6]
  wire  _T_851 = _T_352 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 392307:8]
  wire  _T_854 = _T_350 | _T_851; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 392310:8]
  wire  _T_855 = _T_17 & _T_854; // @[Monitor.scala 147:68 chipyard.TestHarness.SmallBoomConfig.fir 392311:8]
  wire  _T_857 = _T_855 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392313:8]
  wire  _T_858 = ~_T_857; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392314:8]
  wire  _T_877 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 392360:6]
  wire  _T_879 = _T_877 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392362:6]
  wire  _T_880 = ~_T_879; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392363:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.SmallBoomConfig.fir 392368:6]
  wire  _T_881 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 392373:6]
  wire  _T_883 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392376:8]
  wire  _T_884 = ~_T_883; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392377:8]
  wire  _T_885 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 392382:8]
  wire  _T_887 = _T_885 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392384:8]
  wire  _T_888 = ~_T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392385:8]
  wire  _T_889 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.SmallBoomConfig.fir 392390:8]
  wire  _T_891 = _T_889 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392392:8]
  wire  _T_892 = ~_T_891; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392393:8]
  wire  _T_893 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.SmallBoomConfig.fir 392398:8]
  wire  _T_895 = _T_893 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392400:8]
  wire  _T_896 = ~_T_895; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392401:8]
  wire  _T_897 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.SmallBoomConfig.fir 392406:8]
  wire  _T_899 = _T_897 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392408:8]
  wire  _T_900 = ~_T_899; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392409:8]
  wire  _T_901 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 392415:6]
  wire  _T_912 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.SmallBoomConfig.fir 392439:8]
  wire  _T_914 = _T_912 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392441:8]
  wire  _T_915 = ~_T_914; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392442:8]
  wire  _T_916 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.SmallBoomConfig.fir 392447:8]
  wire  _T_918 = _T_916 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392449:8]
  wire  _T_919 = ~_T_918; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392450:8]
  wire  _T_929 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 392473:6]
  wire  _T_949 = _T_897 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.SmallBoomConfig.fir 392514:8]
  wire  _T_951 = _T_949 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392516:8]
  wire  _T_952 = ~_T_951; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392517:8]
  wire  _T_958 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 392532:6]
  wire  _T_975 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 392567:6]
  wire  _T_993 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 392603:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 392669:4]
  wire [8:0] a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 392674:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 392676:4]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392678:4]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 392680:4]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 392681:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 392692:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 392694:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 392696:4]
  wire  _T_1022 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 392697:4]
  wire  _T_1023 = io_in_a_valid & _T_1022; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 392698:4]
  wire  _T_1024 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 392700:6]
  wire  _T_1026 = _T_1024 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392702:6]
  wire  _T_1027 = ~_T_1026; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392703:6]
  wire  _T_1032 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 392716:6]
  wire  _T_1034 = _T_1032 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392718:6]
  wire  _T_1035 = ~_T_1034; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392719:6]
  wire  _T_1040 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 392732:6]
  wire  _T_1042 = _T_1040 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392734:6]
  wire  _T_1043 = ~_T_1042; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392735:6]
  wire  _T_1045 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 392742:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 392750:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 392752:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 392754:4]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 392755:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 392756:4]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392758:4]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 392760:4]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 392761:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 392772:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.SmallBoomConfig.fir 392773:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 392774:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 392775:4]
  reg [2:0] sink; // @[Monitor.scala 539:22 chipyard.TestHarness.SmallBoomConfig.fir 392776:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.SmallBoomConfig.fir 392777:4]
  wire  _T_1046 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 392778:4]
  wire  _T_1047 = io_in_d_valid & _T_1046; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 392779:4]
  wire  _T_1048 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 392781:6]
  wire  _T_1050 = _T_1048 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392783:6]
  wire  _T_1051 = ~_T_1050; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392784:6]
  wire  _T_1052 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.SmallBoomConfig.fir 392789:6]
  wire  _T_1054 = _T_1052 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392791:6]
  wire  _T_1055 = ~_T_1054; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392792:6]
  wire  _T_1056 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 392797:6]
  wire  _T_1058 = _T_1056 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392799:6]
  wire  _T_1059 = ~_T_1058; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392800:6]
  wire  _T_1060 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 392805:6]
  wire  _T_1062 = _T_1060 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392807:6]
  wire  _T_1063 = ~_T_1062; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392808:6]
  wire  _T_1064 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.SmallBoomConfig.fir 392813:6]
  wire  _T_1066 = _T_1064 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392815:6]
  wire  _T_1067 = ~_T_1066; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392816:6]
  wire  _T_1068 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.SmallBoomConfig.fir 392821:6]
  wire  _T_1070 = _T_1068 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392823:6]
  wire  _T_1071 = ~_T_1070; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392824:6]
  wire  _T_1073 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 392831:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 392840:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 392841:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 392842:4]
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392852:4]
  wire [8:0] a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 392854:4]
  wire  a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 392855:4]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392874:4]
  wire [8:0] d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 392876:4]
  wire  d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 392877:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 392898:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 392898:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 392899:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 392903:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 392904:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 392904:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 392905:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.SmallBoomConfig.fir 392909:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 392910:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 392914:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 392915:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 392915:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 392916:4]
  wire  _T_1074 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 392940:4]
  wire [1:0] _GEN_15 = _T_1074 ? 2'h1 : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 392942:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 392944:6 chipyard.TestHarness.SmallBoomConfig.fir 392891:4]
  wire  _T_1077 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 392947:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 392952:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 392953:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 392955:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 392956:6]
  wire [3:0] a_opcodes_set_interm = _T_1077 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392949:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 392954:6 chipyard.TestHarness.SmallBoomConfig.fir 392937:4]
  wire [18:0] _a_opcodes_set_T_1 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 392959:6]
  wire [4:0] a_sizes_set_interm = _T_1077 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392949:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 392957:6 chipyard.TestHarness.SmallBoomConfig.fir 392939:4]
  wire [19:0] _a_sizes_set_T_1 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 392962:6]
  wire  _T_1081 = ~inflight; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 392966:6]
  wire  _T_1083 = _T_1081 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392968:6]
  wire  _T_1084 = ~_T_1083; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392969:6]
  wire [1:0] _GEN_16 = _T_1077 ? 2'h1 : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392949:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 392951:6 chipyard.TestHarness.SmallBoomConfig.fir 392889:4]
  wire [18:0] _GEN_19 = _T_1077 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392949:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 392960:6 chipyard.TestHarness.SmallBoomConfig.fir 392893:4]
  wire [19:0] _GEN_20 = _T_1077 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392949:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 392963:6 chipyard.TestHarness.SmallBoomConfig.fir 392895:4]
  wire  _T_1085 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 392984:4]
  wire  _T_1087 = ~_T_881; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 392986:4]
  wire  _T_1088 = _T_1085 & _T_1087; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 392987:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 392989:6]
  wire [1:0] _GEN_21 = _T_1088 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 392988:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 392990:6 chipyard.TestHarness.SmallBoomConfig.fir 392978:4]
  wire  _T_1090 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 392993:4]
  wire  _T_1093 = _T_1090 & _T_1087; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 392996:4]
  wire [30:0] _GEN_78 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 393005:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_78 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 393005:6]
  wire [30:0] _GEN_79 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.SmallBoomConfig.fir 393012:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_79 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.SmallBoomConfig.fir 393012:6]
  wire [1:0] _GEN_22 = _T_1093 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 392997:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 392999:6 chipyard.TestHarness.SmallBoomConfig.fir 392976:4]
  wire [30:0] _GEN_23 = _T_1093 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 392997:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 393006:6 chipyard.TestHarness.SmallBoomConfig.fir 392980:4]
  wire [30:0] _GEN_24 = _T_1093 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 392997:4 Monitor.scala 678:21 chipyard.TestHarness.SmallBoomConfig.fir 393013:6 chipyard.TestHarness.SmallBoomConfig.fir 392982:4]
  wire  same_cycle_resp = _T_1074 & _source_ok_T_1; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 393023:6]
  wire  _T_1098 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 393024:6]
  wire  _T_1100 = _T_1098 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 393026:6]
  wire  _T_1102 = _T_1100 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393028:6]
  wire  _T_1103 = ~_T_1102; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393029:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8]
  wire  _T_1104 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 393035:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 393036:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 393036:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 393036:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 393036:8]
  wire  _T_1105 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 393036:8]
  wire  _T_1106 = _T_1104 | _T_1105; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 393037:8]
  wire  _T_1108 = _T_1106 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393039:8]
  wire  _T_1109 = ~_T_1108; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393040:8]
  wire  _T_1110 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 393045:8]
  wire  _T_1112 = _T_1110 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393047:8]
  wire  _T_1113 = ~_T_1112; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393048:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392896:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 392906:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8]
  wire  _T_1115 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 393056:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 393058:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 393058:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 393058:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 393058:8]
  wire  _T_1117 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 393058:8]
  wire  _T_1118 = _T_1115 | _T_1117; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 393059:8]
  wire  _T_1120 = _T_1118 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393061:8]
  wire  _T_1121 = ~_T_1120; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393062:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392907:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 392917:4]
  wire [7:0] _GEN_80 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 393067:8]
  wire  _T_1122 = _GEN_80 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 393067:8]
  wire  _T_1124 = _T_1122 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393069:8]
  wire  _T_1125 = ~_T_1124; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393070:8]
  wire  _T_1127 = _T_1085 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 393078:4]
  wire  _T_1128 = _T_1127 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 393079:4]
  wire  _T_1130 = _T_1128 & _source_ok_T_1; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 393081:4]
  wire  _T_1132 = _T_1130 & _T_1087; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 393083:4]
  wire  _T_1133 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 393085:6]
  wire  _T_1134 = _T_1133 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 393086:6]
  wire  _T_1136 = _T_1134 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393088:6]
  wire  _T_1137 = ~_T_1136; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393089:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392890:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392977:4]
  wire  _T_1138 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 393095:4]
  wire  _T_1139 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 393096:4]
  wire  _T_1140 = ~_T_1139; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 393097:4]
  wire  _T_1141 = _T_1138 | _T_1140; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 393098:4]
  wire  _T_1143 = _T_1141 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393100:4]
  wire  _T_1144 = ~_T_1143; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393101:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392888:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 393106:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392975:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 393107:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 393108:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392892:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 393110:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392979:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 393111:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 393112:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392894:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 393114:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392981:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.SmallBoomConfig.fir 393115:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 393116:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 393118:4]
  wire  _T_1145 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 393121:4]
  wire  _T_1146 = ~_T_1145; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 393122:4]
  wire  _T_1147 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 393123:4]
  wire  _T_1148 = _T_1146 | _T_1147; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 393124:4]
  wire  _T_1149 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 393125:4]
  wire  _T_1150 = _T_1148 | _T_1149; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 393126:4]
  wire  _T_1152 = _T_1150 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 393128:4]
  wire  _T_1153 = ~_T_1152; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 393129:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 393135:4]
  wire  _T_1156 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 393139:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 393145:4]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 393180:4]
  wire [8:0] d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 393182:4]
  wire  d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 393183:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 393216:4]
  wire [15:0] _GEN_84 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 393221:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_84 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 393221:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 393222:4]
  wire  _T_1174 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 393300:4]
  wire  _T_1176 = _T_1174 & _T_881; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 393302:4]
  wire  _T_1178 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 393308:4]
  wire  _T_1180 = _T_1178 & _T_881; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 393310:4]
  wire [30:0] _GEN_69 = _T_1180 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 393311:4 Monitor.scala 786:21 chipyard.TestHarness.SmallBoomConfig.fir 393327:6 chipyard.TestHarness.SmallBoomConfig.fir 393298:4]
  wire  _T_1184 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 393346:6]
  wire  _T_1188 = _T_1184 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393350:6]
  wire  _T_1189 = ~_T_1188; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393351:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 393204:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 393223:4]
  wire  _T_1194 = _GEN_80 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 393369:8]
  wire  _T_1196 = _T_1194 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393371:8]
  wire  _T_1197 = ~_T_1196; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393372:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 393297:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.SmallBoomConfig.fir 393422:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 393423:4]
  wire  _GEN_90 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391352:10]
  wire  _GEN_100 = io_in_a_valid & _T_171; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391542:10]
  wire  _GEN_112 = io_in_a_valid & _T_331; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391680:10]
  wire  _GEN_120 = io_in_a_valid & _T_426; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391872:10]
  wire  _GEN_126 = io_in_a_valid & _T_517; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391985:10]
  wire  _GEN_132 = io_in_a_valid & _T_610; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392095:10]
  wire  _GEN_138 = io_in_a_valid & _T_696; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392203:10]
  wire  _GEN_144 = io_in_a_valid & _T_782; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392316:10]
  wire  _GEN_150 = io_in_d_valid & _T_881; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392379:10]
  wire  _GEN_160 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392421:10]
  wire  _GEN_170 = io_in_d_valid & _T_929; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392479:10]
  wire  _GEN_180 = io_in_d_valid & _T_958; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392538:10]
  wire  _GEN_186 = io_in_d_valid & _T_975; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392573:10]
  wire  _GEN_192 = io_in_d_valid & _T_993; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392609:10]
  wire  _GEN_198 = _T_1088 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393042:10]
  wire  _GEN_203 = _T_1088 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393064:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 393119:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 393426:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392678:4]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392678:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 392688:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 392689:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392677:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 392743:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 392744:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 392743:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 392746:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 392743:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 392748:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392758:4]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392758:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 392768:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 392769:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392757:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392832:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 392833:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392832:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.SmallBoomConfig.fir 392834:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392832:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 392835:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392832:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 392836:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392832:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.SmallBoomConfig.fir 392837:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392832:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.SmallBoomConfig.fir 392838:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 392840:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 392840:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 393109:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 392841:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 392841:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 393113:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 392842:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 392842:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 393117:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392852:4]
      a_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392852:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 392862:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 392863:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392677:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392874:4]
      d_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392874:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 392884:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 392885:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392757:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 393118:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 393118:4]
    end else if (_T_1156) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 393140:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 393141:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 393136:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 393145:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 393145:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 393424:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 393180:4]
      d_first_counter_2 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 393180:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 393190:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 393191:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392757:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391352:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391353:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391419:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391420:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391434:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391435:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391441:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391442:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391458:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391459:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391542:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391543:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391609:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391610:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391624:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391625:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391631:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391632:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391647:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391648:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391656:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391657:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_331 & _T_340) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391680:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_340) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391681:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_407) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391751:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_407) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391752:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391765:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391766:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391781:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391782:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_426 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391872:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391873:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391886:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391887:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391902:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391903:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_517 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391985:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391986:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391999:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392000:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392017:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392018:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_610 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392095:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392096:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392109:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392110:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392125:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392126:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_696 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392203:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392204:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392217:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392218:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392233:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392234:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_782 & _T_858) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392316:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_858) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392317:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392330:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392331:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392346:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392347:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392365:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392366:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_881 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392379:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392380:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392387:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392388:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392395:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392396:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392403:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392404:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_900) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392411:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_900) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392412:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_901 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392421:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392422:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392436:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392437:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392444:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392445:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392452:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392453:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392460:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392461:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_929 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392479:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392480:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392494:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392495:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392502:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392503:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392510:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392511:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392519:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392520:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_958 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392538:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392539:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392546:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392547:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392554:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392555:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_975 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392573:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392574:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392581:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392582:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392590:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392591:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_993 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392609:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392610:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392617:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392618:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392625:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392626:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392705:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392706:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392721:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392722:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392737:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392738:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392786:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392787:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392794:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392795:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392802:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392803:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392810:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392811:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392818:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392819:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392826:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392827:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392971:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392972:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393031:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393032:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & same_cycle_resp & _T_1109) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393042:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_1109) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393043:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_1113) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393050:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_1113) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393051:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & ~same_cycle_resp & _T_1121) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393064:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_1121) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393065:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_1125) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393072:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_1125) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393073:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393091:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393092:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1144) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 8 (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393103:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1144) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393104:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1153) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 393131:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1153) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 393132:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393353:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393354:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393374:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393375:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  address = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  d_first_counter = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  opcode_1 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  param_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  size_1 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  source_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sink = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  denied = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inflight = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight_opcodes = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  inflight_sizes = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  watchdog = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_21_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393581:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393582:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393583:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [3:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [31:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output        auto_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [3:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input         auto_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [2:0]  auto_out_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire [2:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire  bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  TLMonitor_57_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393591:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_6_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393618:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_7_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 393630:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393631:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 393644:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393592:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393593:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 393630:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393619:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393620:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393633:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393614:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393616:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393589:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393617:4]
endmodule
module SerialRAM_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393665:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393666:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393667:4]
  input         io_ser_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  output        io_ser_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  output [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  output        io_ser_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  input         io_ser_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  input  [3:0]  io_ser_out_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  output        io_tsi_ser_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  input         io_tsi_ser_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  input  [31:0] io_tsi_ser_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  input         io_tsi_ser_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  output        io_tsi_ser_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  output [31:0] io_tsi_ser_out_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
);
  wire  adapter_clock; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_reset; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_auto_out_a_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_auto_out_a_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire [2:0] adapter_auto_out_a_bits_opcode; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire [3:0] adapter_auto_out_a_bits_size; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire [31:0] adapter_auto_out_a_bits_address; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire [7:0] adapter_auto_out_a_bits_mask; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire [63:0] adapter_auto_out_a_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_auto_out_d_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_auto_out_d_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire [63:0] adapter_auto_out_d_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_io_serial_in_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_io_serial_in_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire [31:0] adapter_io_serial_in_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_io_serial_out_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  adapter_io_serial_out_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire [31:0] adapter_io_serial_out_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  wire  serdesser_clock; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_reset; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [3:0] serdesser_auto_manager_in_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [31:0] serdesser_auto_manager_in_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [7:0] serdesser_auto_manager_in_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [63:0] serdesser_auto_manager_in_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [1:0] serdesser_auto_manager_in_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [3:0] serdesser_auto_manager_in_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [63:0] serdesser_auto_manager_in_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_manager_in_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_client_out_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_client_out_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_client_out_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_client_out_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_client_out_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [3:0] serdesser_auto_client_out_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [28:0] serdesser_auto_client_out_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [7:0] serdesser_auto_client_out_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [63:0] serdesser_auto_client_out_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_client_out_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_client_out_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_client_out_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_client_out_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [1:0] serdesser_auto_client_out_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [2:0] serdesser_auto_client_out_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [3:0] serdesser_auto_client_out_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_client_out_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_client_out_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [63:0] serdesser_auto_client_out_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_auto_client_out_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_io_ser_in_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_io_ser_in_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [3:0] serdesser_io_ser_in_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_io_ser_out_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  serdesser_io_ser_out_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire [3:0] serdesser_io_ser_out_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
  wire  srams_clock; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire  srams_reset; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire  srams_auto_in_a_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire  srams_auto_in_a_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [2:0] srams_auto_in_a_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [2:0] srams_auto_in_a_bits_param; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [1:0] srams_auto_in_a_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [7:0] srams_auto_in_a_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [28:0] srams_auto_in_a_bits_address; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [7:0] srams_auto_in_a_bits_mask; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [63:0] srams_auto_in_a_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire  srams_auto_in_a_bits_corrupt; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire  srams_auto_in_d_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire  srams_auto_in_d_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [2:0] srams_auto_in_d_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [1:0] srams_auto_in_d_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [7:0] srams_auto_in_d_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire [63:0] srams_auto_in_d_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
  wire  xbar_auto_in_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_in_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_in_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_in_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_in_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [3:0] xbar_auto_in_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [28:0] xbar_auto_in_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [7:0] xbar_auto_in_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [63:0] xbar_auto_in_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_in_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_in_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_in_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_in_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [1:0] xbar_auto_in_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_in_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [3:0] xbar_auto_in_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_in_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_in_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [63:0] xbar_auto_in_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_in_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_out_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_out_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_out_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_out_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_out_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [3:0] xbar_auto_out_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [28:0] xbar_auto_out_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [7:0] xbar_auto_out_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [63:0] xbar_auto_out_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_out_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_out_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_out_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_out_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [1:0] xbar_auto_out_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [2:0] xbar_auto_out_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [3:0] xbar_auto_out_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_out_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_out_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire [63:0] xbar_auto_out_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  xbar_auto_out_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
  wire  buffer_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [1:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [7:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [28:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_in_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [1:0] buffer_auto_in_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [1:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [7:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_in_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [1:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [7:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [28:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [1:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [7:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [2:0] fragmenter_auto_in_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [3:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [28:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [63:0] fragmenter_auto_in_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_in_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [1:0] fragmenter_auto_in_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [3:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_in_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_in_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_in_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [2:0] fragmenter_auto_out_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [7:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [28:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [7:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [63:0] fragmenter_auto_out_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_out_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [1:0] fragmenter_auto_out_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [7:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_out_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_out_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  fragmenter_auto_out_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  buffer_1_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [2:0] buffer_1_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [3:0] buffer_1_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [31:0] buffer_1_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [7:0] buffer_1_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [63:0] buffer_1_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [63:0] buffer_1_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [2:0] buffer_1_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [2:0] buffer_1_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [3:0] buffer_1_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [31:0] buffer_1_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [7:0] buffer_1_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [63:0] buffer_1_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [2:0] buffer_1_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [1:0] buffer_1_auto_out_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [3:0] buffer_1_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [2:0] buffer_1_auto_out_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire [63:0] buffer_1_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  wire  buffer_1_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
  SerialAdapter_inTestHarness adapter ( // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
    .clock(adapter_clock),
    .reset(adapter_reset),
    .auto_out_a_ready(adapter_auto_out_a_ready),
    .auto_out_a_valid(adapter_auto_out_a_valid),
    .auto_out_a_bits_opcode(adapter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(adapter_auto_out_a_bits_size),
    .auto_out_a_bits_address(adapter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(adapter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(adapter_auto_out_a_bits_data),
    .auto_out_d_ready(adapter_auto_out_d_ready),
    .auto_out_d_valid(adapter_auto_out_d_valid),
    .auto_out_d_bits_data(adapter_auto_out_d_bits_data),
    .io_serial_in_ready(adapter_io_serial_in_ready),
    .io_serial_in_valid(adapter_io_serial_in_valid),
    .io_serial_in_bits(adapter_io_serial_in_bits),
    .io_serial_out_ready(adapter_io_serial_out_ready),
    .io_serial_out_valid(adapter_io_serial_out_valid),
    .io_serial_out_bits(adapter_io_serial_out_bits)
  );
  TLSerdesser_1_inTestHarness serdesser ( // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393682:4]
    .clock(serdesser_clock),
    .reset(serdesser_reset),
    .auto_manager_in_a_ready(serdesser_auto_manager_in_a_ready),
    .auto_manager_in_a_valid(serdesser_auto_manager_in_a_valid),
    .auto_manager_in_a_bits_opcode(serdesser_auto_manager_in_a_bits_opcode),
    .auto_manager_in_a_bits_param(serdesser_auto_manager_in_a_bits_param),
    .auto_manager_in_a_bits_size(serdesser_auto_manager_in_a_bits_size),
    .auto_manager_in_a_bits_source(serdesser_auto_manager_in_a_bits_source),
    .auto_manager_in_a_bits_address(serdesser_auto_manager_in_a_bits_address),
    .auto_manager_in_a_bits_mask(serdesser_auto_manager_in_a_bits_mask),
    .auto_manager_in_a_bits_data(serdesser_auto_manager_in_a_bits_data),
    .auto_manager_in_a_bits_corrupt(serdesser_auto_manager_in_a_bits_corrupt),
    .auto_manager_in_d_ready(serdesser_auto_manager_in_d_ready),
    .auto_manager_in_d_valid(serdesser_auto_manager_in_d_valid),
    .auto_manager_in_d_bits_opcode(serdesser_auto_manager_in_d_bits_opcode),
    .auto_manager_in_d_bits_param(serdesser_auto_manager_in_d_bits_param),
    .auto_manager_in_d_bits_size(serdesser_auto_manager_in_d_bits_size),
    .auto_manager_in_d_bits_source(serdesser_auto_manager_in_d_bits_source),
    .auto_manager_in_d_bits_sink(serdesser_auto_manager_in_d_bits_sink),
    .auto_manager_in_d_bits_denied(serdesser_auto_manager_in_d_bits_denied),
    .auto_manager_in_d_bits_data(serdesser_auto_manager_in_d_bits_data),
    .auto_manager_in_d_bits_corrupt(serdesser_auto_manager_in_d_bits_corrupt),
    .auto_client_out_a_ready(serdesser_auto_client_out_a_ready),
    .auto_client_out_a_valid(serdesser_auto_client_out_a_valid),
    .auto_client_out_a_bits_opcode(serdesser_auto_client_out_a_bits_opcode),
    .auto_client_out_a_bits_param(serdesser_auto_client_out_a_bits_param),
    .auto_client_out_a_bits_size(serdesser_auto_client_out_a_bits_size),
    .auto_client_out_a_bits_source(serdesser_auto_client_out_a_bits_source),
    .auto_client_out_a_bits_address(serdesser_auto_client_out_a_bits_address),
    .auto_client_out_a_bits_mask(serdesser_auto_client_out_a_bits_mask),
    .auto_client_out_a_bits_data(serdesser_auto_client_out_a_bits_data),
    .auto_client_out_a_bits_corrupt(serdesser_auto_client_out_a_bits_corrupt),
    .auto_client_out_d_ready(serdesser_auto_client_out_d_ready),
    .auto_client_out_d_valid(serdesser_auto_client_out_d_valid),
    .auto_client_out_d_bits_opcode(serdesser_auto_client_out_d_bits_opcode),
    .auto_client_out_d_bits_param(serdesser_auto_client_out_d_bits_param),
    .auto_client_out_d_bits_size(serdesser_auto_client_out_d_bits_size),
    .auto_client_out_d_bits_source(serdesser_auto_client_out_d_bits_source),
    .auto_client_out_d_bits_sink(serdesser_auto_client_out_d_bits_sink),
    .auto_client_out_d_bits_denied(serdesser_auto_client_out_d_bits_denied),
    .auto_client_out_d_bits_data(serdesser_auto_client_out_d_bits_data),
    .auto_client_out_d_bits_corrupt(serdesser_auto_client_out_d_bits_corrupt),
    .io_ser_in_ready(serdesser_io_ser_in_ready),
    .io_ser_in_valid(serdesser_io_ser_in_valid),
    .io_ser_in_bits(serdesser_io_ser_in_bits),
    .io_ser_out_ready(serdesser_io_ser_out_ready),
    .io_ser_out_valid(serdesser_io_ser_out_valid),
    .io_ser_out_bits(serdesser_io_ser_out_bits)
  );
  TLRAM_inTestHarness srams ( // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393689:4]
    .clock(srams_clock),
    .reset(srams_reset),
    .auto_in_a_ready(srams_auto_in_a_ready),
    .auto_in_a_valid(srams_auto_in_a_valid),
    .auto_in_a_bits_opcode(srams_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(srams_auto_in_a_bits_param),
    .auto_in_a_bits_size(srams_auto_in_a_bits_size),
    .auto_in_a_bits_source(srams_auto_in_a_bits_source),
    .auto_in_a_bits_address(srams_auto_in_a_bits_address),
    .auto_in_a_bits_mask(srams_auto_in_a_bits_mask),
    .auto_in_a_bits_data(srams_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(srams_auto_in_a_bits_corrupt),
    .auto_in_d_ready(srams_auto_in_d_ready),
    .auto_in_d_valid(srams_auto_in_d_valid),
    .auto_in_d_bits_opcode(srams_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(srams_auto_in_d_bits_size),
    .auto_in_d_bits_source(srams_auto_in_d_bits_source),
    .auto_in_d_bits_data(srams_auto_in_d_bits_data)
  );
  TLXbar_10_inTestHarness xbar ( // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393695:4]
    .auto_in_a_ready(xbar_auto_in_a_ready),
    .auto_in_a_valid(xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(xbar_auto_in_a_bits_corrupt),
    .auto_in_d_ready(xbar_auto_in_d_ready),
    .auto_in_d_valid(xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(xbar_auto_out_a_ready),
    .auto_out_a_valid(xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(xbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(xbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(xbar_auto_out_a_bits_corrupt),
    .auto_out_d_ready(xbar_auto_out_d_ready),
    .auto_out_d_valid(xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(xbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(xbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(xbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(xbar_auto_out_d_bits_corrupt)
  );
  TLBuffer_20_inTestHarness buffer ( // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data)
  );
  TLFragmenter_7_inTestHarness fragmenter ( // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fragmenter_auto_in_d_bits_param),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fragmenter_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fragmenter_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fragmenter_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fragmenter_auto_out_d_bits_param),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fragmenter_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fragmenter_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fragmenter_auto_out_d_bits_corrupt)
  );
  TLBuffer_21_inTestHarness buffer_1 ( // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393713:4]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_a_ready(buffer_1_auto_in_a_ready),
    .auto_in_a_valid(buffer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
    .auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_1_auto_in_d_ready),
    .auto_in_d_valid(buffer_1_auto_in_d_valid),
    .auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
    .auto_out_a_ready(buffer_1_auto_out_a_ready),
    .auto_out_a_valid(buffer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_1_auto_out_d_ready),
    .auto_out_d_valid(buffer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
  );
  assign io_ser_in_valid = serdesser_io_ser_out_valid; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.SmallBoomConfig.fir 393729:4]
  assign io_ser_in_bits = serdesser_io_ser_out_bits; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.SmallBoomConfig.fir 393728:4]
  assign io_ser_out_ready = serdesser_io_ser_in_ready; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.SmallBoomConfig.fir 393727:4]
  assign io_tsi_ser_in_ready = adapter_io_serial_in_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393736:4]
  assign io_tsi_ser_out_valid = adapter_io_serial_out_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393732:4]
  assign io_tsi_ser_out_bits = adapter_io_serial_out_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393731:4]
  assign adapter_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393680:4]
  assign adapter_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393681:4]
  assign adapter_auto_out_a_ready = buffer_1_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign adapter_auto_out_d_valid = buffer_1_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign adapter_auto_out_d_bits_data = buffer_1_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign adapter_io_serial_in_valid = io_tsi_ser_in_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393735:4]
  assign adapter_io_serial_in_bits = io_tsi_ser_in_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393734:4]
  assign adapter_io_serial_out_ready = io_tsi_ser_out_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393733:4]
  assign serdesser_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393687:4]
  assign serdesser_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393688:4]
  assign serdesser_auto_manager_in_a_valid = buffer_1_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_a_bits_param = buffer_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_a_bits_size = buffer_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_a_bits_source = buffer_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_a_bits_address = buffer_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_a_bits_data = buffer_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_manager_in_d_ready = buffer_1_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign serdesser_auto_client_out_a_ready = xbar_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_valid = xbar_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_bits_opcode = xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_bits_param = xbar_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_bits_size = xbar_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_bits_source = xbar_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_bits_sink = xbar_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_bits_denied = xbar_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_bits_data = xbar_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_auto_client_out_d_bits_corrupt = xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign serdesser_io_ser_in_valid = io_ser_out_valid; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.SmallBoomConfig.fir 393726:4]
  assign serdesser_io_ser_in_bits = io_ser_out_bits; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.SmallBoomConfig.fir 393725:4]
  assign serdesser_io_ser_out_ready = io_ser_in_ready; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.SmallBoomConfig.fir 393730:4]
  assign srams_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393693:4]
  assign srams_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393694:4]
  assign srams_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign srams_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign xbar_auto_in_a_valid = serdesser_auto_client_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_a_bits_opcode = serdesser_auto_client_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_a_bits_param = serdesser_auto_client_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_a_bits_size = serdesser_auto_client_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_a_bits_source = serdesser_auto_client_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_a_bits_address = serdesser_auto_client_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_a_bits_mask = serdesser_auto_client_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_a_bits_data = serdesser_auto_client_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_a_bits_corrupt = serdesser_auto_client_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_in_d_ready = serdesser_auto_client_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393720:4]
  assign xbar_auto_out_a_ready = fragmenter_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_valid = fragmenter_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_bits_param = fragmenter_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_bits_sink = fragmenter_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_bits_denied = fragmenter_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign xbar_auto_out_d_bits_corrupt = fragmenter_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign buffer_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393705:4]
  assign buffer_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393706:4]
  assign buffer_auto_in_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_a_bits_param = fragmenter_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_a_bits_data = fragmenter_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_in_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_auto_out_a_ready = srams_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign buffer_auto_out_d_valid = srams_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign buffer_auto_out_d_bits_opcode = srams_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign buffer_auto_out_d_bits_size = srams_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign buffer_auto_out_d_bits_source = srams_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign buffer_auto_out_d_bits_data = srams_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393722:4]
  assign fragmenter_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393711:4]
  assign fragmenter_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393712:4]
  assign fragmenter_auto_in_a_valid = xbar_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_a_bits_opcode = xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_a_bits_param = xbar_auto_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_a_bits_size = xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_a_bits_source = xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_a_bits_address = xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_a_bits_mask = xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_a_bits_data = xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_a_bits_corrupt = xbar_auto_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_in_d_ready = xbar_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393721:4]
  assign fragmenter_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign fragmenter_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393723:4]
  assign buffer_1_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393717:4]
  assign buffer_1_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393718:4]
  assign buffer_1_auto_in_a_valid = adapter_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign buffer_1_auto_in_a_bits_opcode = adapter_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign buffer_1_auto_in_a_bits_size = adapter_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign buffer_1_auto_in_a_bits_address = adapter_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign buffer_1_auto_in_a_bits_mask = adapter_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign buffer_1_auto_in_a_bits_data = adapter_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign buffer_1_auto_in_d_ready = adapter_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393719:4]
  assign buffer_1_auto_out_a_ready = serdesser_auto_manager_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_valid = serdesser_auto_manager_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_bits_opcode = serdesser_auto_manager_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_bits_param = serdesser_auto_manager_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_bits_size = serdesser_auto_manager_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_bits_source = serdesser_auto_manager_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_bits_sink = serdesser_auto_manager_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_bits_denied = serdesser_auto_manager_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_bits_data = serdesser_auto_manager_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
  assign buffer_1_auto_out_d_bits_corrupt = serdesser_auto_manager_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393724:4]
endmodule
module Queue_48_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393759:2]
  input        clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393760:4]
  input        reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393761:4]
  output       io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393762:4]
  input        io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393762:4]
  input  [7:0] io_enq_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 393762:4]
  input        io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393762:4]
  output       io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393762:4]
  output [7:0] io_deq_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 393762:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:127]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
  wire [6:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
  wire [6:0] ram_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
  reg [6:0] enq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393765:4]
  reg [6:0] deq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393766:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 393767:4]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 393768:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 393769:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 393770:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 393771:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 393772:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 393775:4]
  wire [6:0] _value_T_1 = enq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393783:6]
  wire [6:0] _value_T_3 = deq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393789:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 393792:4]
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 393798:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 393796:4]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 393801:4]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393764:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393765:4]
      enq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393765:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 393778:4]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393784:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393766:4]
      deq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393766:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 393786:4]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393790:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 393767:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 393767:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 393793:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 393794:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UARTAdapter_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393867:2]
  input   clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393868:4]
  input   reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393869:4]
  input   io_uart_txd, // @[chipyard.TestHarness.SmallBoomConfig.fir 393870:4]
  output  io_uart_rxd // @[chipyard.TestHarness.SmallBoomConfig.fir 393870:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  txfifo_clock; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
  wire  txfifo_reset; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
  wire  txfifo_io_enq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
  wire  txfifo_io_enq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
  wire [7:0] txfifo_io_enq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
  wire  txfifo_io_deq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
  wire  txfifo_io_deq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
  wire [7:0] txfifo_io_deq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
  wire  rxfifo_clock; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
  wire  rxfifo_reset; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
  wire  rxfifo_io_enq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
  wire  rxfifo_io_enq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
  wire [7:0] rxfifo_io_enq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
  wire  rxfifo_io_deq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
  wire  rxfifo_io_deq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
  wire [7:0] rxfifo_io_deq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
  wire  sim_clock; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
  wire  sim_reset; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
  wire  sim_serial_in_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
  wire  sim_serial_in_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
  wire [7:0] sim_serial_in_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
  wire  sim_serial_out_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
  wire  sim_serial_out_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
  wire [7:0] sim_serial_out_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
  reg [1:0] txState; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393878:4]
  reg [7:0] txData; // @[UARTAdapter.scala 39:19 chipyard.TestHarness.SmallBoomConfig.fir 393879:4]
  wire  _T = txState == 2'h2; // @[UARTAdapter.scala 41:49 chipyard.TestHarness.SmallBoomConfig.fir 393880:4]
  wire  _T_1 = _T & txfifo_io_enq_ready; // @[UARTAdapter.scala 41:61 chipyard.TestHarness.SmallBoomConfig.fir 393881:4]
  reg [2:0] txDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393882:4]
  wire  wrap_wrap = txDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393886:6]
  wire [2:0] _wrap_value_T_1 = txDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393888:6]
  wire  txDataWrap = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393885:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393890:6 chipyard.TestHarness.SmallBoomConfig.fir 393884:4]
  wire  _T_2 = txState == 2'h1; // @[UARTAdapter.scala 43:51 chipyard.TestHarness.SmallBoomConfig.fir 393892:4]
  wire  _T_3 = _T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 43:63 chipyard.TestHarness.SmallBoomConfig.fir 393893:4]
  reg [9:0] txBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393894:4]
  wire  wrap_wrap_1 = txBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393898:6]
  wire [9:0] _wrap_value_T_3 = txBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393900:6]
  wire  txBaudWrap = _T_3 & wrap_wrap_1; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393897:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393905:6 chipyard.TestHarness.SmallBoomConfig.fir 393896:4]
  wire  _T_4 = txState == 2'h0; // @[UARTAdapter.scala 44:53 chipyard.TestHarness.SmallBoomConfig.fir 393907:4]
  wire  _T_5 = ~io_uart_txd; // @[UARTAdapter.scala 44:80 chipyard.TestHarness.SmallBoomConfig.fir 393908:4]
  wire  _T_6 = _T_4 & _T_5; // @[UARTAdapter.scala 44:65 chipyard.TestHarness.SmallBoomConfig.fir 393909:4]
  wire  _T_7 = _T_6 & txfifo_io_enq_ready; // @[UARTAdapter.scala 44:88 chipyard.TestHarness.SmallBoomConfig.fir 393910:4]
  reg [1:0] txSlackCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393911:4]
  wire  wrap_wrap_2 = txSlackCount == 2'h3; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393915:6]
  wire [1:0] _wrap_value_T_5 = txSlackCount + 2'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393917:6]
  wire  txSlackWrap = _T_7 & wrap_wrap_2; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393914:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393919:6 chipyard.TestHarness.SmallBoomConfig.fir 393913:4]
  wire  _T_8 = 2'h0 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393921:4]
  wire  _T_9 = 2'h1 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393929:6]
  wire  _T_10 = 2'h2 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393936:8]
  wire [7:0] _GEN_35 = {{7'd0}, io_uart_txd}; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.SmallBoomConfig.fir 393939:12]
  wire [7:0] _txData_T = _GEN_35 << txDataIdx; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.SmallBoomConfig.fir 393939:12]
  wire [7:0] _txData_T_1 = txData | _txData_T; // @[UARTAdapter.scala 60:26 chipyard.TestHarness.SmallBoomConfig.fir 393940:12]
  wire [1:0] _txState_T_1 = io_uart_txd ? 2'h0 : 2'h3; // @[UARTAdapter.scala 63:23 chipyard.TestHarness.SmallBoomConfig.fir 393945:12]
  wire [1:0] _GEN_11 = txfifo_io_enq_ready ? 2'h1 : txState; // @[UARTAdapter.scala 64:39 chipyard.TestHarness.SmallBoomConfig.fir 393949:12 UARTAdapter.scala 65:17 chipyard.TestHarness.SmallBoomConfig.fir 393950:14 UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393878:4]
  wire [1:0] _GEN_12 = txDataWrap ? _txState_T_1 : _GEN_11; // @[UARTAdapter.scala 62:24 chipyard.TestHarness.SmallBoomConfig.fir 393943:10 UARTAdapter.scala 63:17 chipyard.TestHarness.SmallBoomConfig.fir 393946:12]
  wire  _T_11 = 2'h3 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393954:10]
  wire  _T_13 = io_uart_txd & txfifo_io_enq_ready; // @[UARTAdapter.scala 69:32 chipyard.TestHarness.SmallBoomConfig.fir 393957:12]
  wire [1:0] _GEN_13 = _T_13 ? 2'h0 : txState; // @[UARTAdapter.scala 69:56 chipyard.TestHarness.SmallBoomConfig.fir 393958:12 UARTAdapter.scala 70:17 chipyard.TestHarness.SmallBoomConfig.fir 393959:14 UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393878:4]
  wire [1:0] _GEN_14 = _T_11 ? _GEN_13 : txState; // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393955:10 UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393878:4]
  reg [1:0] rxState; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.SmallBoomConfig.fir 393964:4]
  reg [9:0] rxBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393965:4]
  wire  wrap_wrap_3 = rxBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393969:6]
  wire [9:0] _wrap_value_T_7 = rxBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393971:6]
  wire  rxBaudWrap = txfifo_io_enq_ready & wrap_wrap_3; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393968:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393976:6 chipyard.TestHarness.SmallBoomConfig.fir 393967:4]
  wire  _T_14 = rxState == 2'h2; // @[UARTAdapter.scala 83:49 chipyard.TestHarness.SmallBoomConfig.fir 393978:4]
  wire  _T_15 = _T_14 & txfifo_io_enq_ready; // @[UARTAdapter.scala 83:61 chipyard.TestHarness.SmallBoomConfig.fir 393979:4]
  wire  _T_16 = _T_15 & rxBaudWrap; // @[UARTAdapter.scala 83:84 chipyard.TestHarness.SmallBoomConfig.fir 393980:4]
  reg [2:0] rxDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393981:4]
  wire  wrap_wrap_4 = rxDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393985:6]
  wire [2:0] _wrap_value_T_9 = rxDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393987:6]
  wire  rxDataWrap = _T_16 & wrap_wrap_4; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393984:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393989:6 chipyard.TestHarness.SmallBoomConfig.fir 393983:4]
  wire  _T_17 = 2'h0 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393992:4]
  wire  _T_18 = rxBaudWrap & rxfifo_io_deq_valid; // @[UARTAdapter.scala 89:24 chipyard.TestHarness.SmallBoomConfig.fir 393995:6]
  wire  _T_19 = 2'h1 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 394001:6]
  wire  _T_20 = 2'h2 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 394009:8]
  wire [7:0] _io_uart_rxd_T = rxfifo_io_deq_bits >> rxDataIdx; // @[UARTAdapter.scala 100:42 chipyard.TestHarness.SmallBoomConfig.fir 394011:10]
  wire  _T_21 = rxDataWrap & rxBaudWrap; // @[UARTAdapter.scala 101:23 chipyard.TestHarness.SmallBoomConfig.fir 394014:10]
  wire [1:0] _GEN_28 = _T_21 ? 2'h0 : rxState; // @[UARTAdapter.scala 101:38 chipyard.TestHarness.SmallBoomConfig.fir 394015:10 UARTAdapter.scala 102:17 chipyard.TestHarness.SmallBoomConfig.fir 394016:12 UARTAdapter.scala 79:24 chipyard.TestHarness.SmallBoomConfig.fir 393964:4]
  wire  _GEN_29 = _T_20 ? _io_uart_rxd_T[0] : 1'h1; // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 394010:8 UARTAdapter.scala 100:19 chipyard.TestHarness.SmallBoomConfig.fir 394013:10 UARTAdapter.scala 85:15 chipyard.TestHarness.SmallBoomConfig.fir 393991:4]
  wire  _GEN_31 = _T_19 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 394002:6 UARTAdapter.scala 94:19 chipyard.TestHarness.SmallBoomConfig.fir 394003:8]
  wire  _rxfifo_io_deq_ready_T_1 = _T_14 & rxDataWrap; // @[UARTAdapter.scala 106:48 chipyard.TestHarness.SmallBoomConfig.fir 394020:4]
  wire  _rxfifo_io_deq_ready_T_2 = _rxfifo_io_deq_ready_T_1 & rxBaudWrap; // @[UARTAdapter.scala 106:62 chipyard.TestHarness.SmallBoomConfig.fir 394021:4]
  Queue_48_inTestHarness txfifo ( // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393872:4]
    .clock(txfifo_clock),
    .reset(txfifo_reset),
    .io_enq_ready(txfifo_io_enq_ready),
    .io_enq_valid(txfifo_io_enq_valid),
    .io_enq_bits(txfifo_io_enq_bits),
    .io_deq_ready(txfifo_io_deq_ready),
    .io_deq_valid(txfifo_io_deq_valid),
    .io_deq_bits(txfifo_io_deq_bits)
  );
  Queue_48_inTestHarness rxfifo ( // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393875:4]
    .clock(rxfifo_clock),
    .reset(rxfifo_reset),
    .io_enq_ready(rxfifo_io_enq_ready),
    .io_enq_valid(rxfifo_io_enq_valid),
    .io_enq_bits(rxfifo_io_enq_bits),
    .io_deq_ready(rxfifo_io_deq_ready),
    .io_deq_valid(rxfifo_io_deq_valid),
    .io_deq_bits(rxfifo_io_deq_bits)
  );
  SimUART #(.UARTNO(0)) sim ( // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 394024:4]
    .clock(sim_clock),
    .reset(sim_reset),
    .serial_in_ready(sim_serial_in_ready),
    .serial_in_valid(sim_serial_in_valid),
    .serial_in_bits(sim_serial_in_bits),
    .serial_out_ready(sim_serial_out_ready),
    .serial_out_valid(sim_serial_out_valid),
    .serial_out_bits(sim_serial_out_bits)
  );
  assign io_uart_rxd = _T_17 | _GEN_31; // @[Conditional.scala 40:58 chipyard.TestHarness.SmallBoomConfig.fir 393993:4 UARTAdapter.scala 88:19 chipyard.TestHarness.SmallBoomConfig.fir 393994:6]
  assign txfifo_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393873:4]
  assign txfifo_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393874:4]
  assign txfifo_io_enq_valid = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393885:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393890:6 chipyard.TestHarness.SmallBoomConfig.fir 393884:4]
  assign txfifo_io_enq_bits = txData; // @[UARTAdapter.scala 75:23 chipyard.TestHarness.SmallBoomConfig.fir 393962:4]
  assign txfifo_io_deq_ready = sim_serial_out_ready; // @[UARTAdapter.scala 115:23 chipyard.TestHarness.SmallBoomConfig.fir 394033:4]
  assign rxfifo_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393876:4]
  assign rxfifo_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393877:4]
  assign rxfifo_io_enq_valid = sim_serial_in_valid; // @[UARTAdapter.scala 118:23 chipyard.TestHarness.SmallBoomConfig.fir 394035:4]
  assign rxfifo_io_enq_bits = sim_serial_in_bits; // @[UARTAdapter.scala 117:22 chipyard.TestHarness.SmallBoomConfig.fir 394034:4]
  assign rxfifo_io_deq_ready = _rxfifo_io_deq_ready_T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 106:76 chipyard.TestHarness.SmallBoomConfig.fir 394022:4]
  assign sim_clock = clock; // @[UARTAdapter.scala 110:16 chipyard.TestHarness.SmallBoomConfig.fir 394028:4]
  assign sim_reset = reset; // @[UARTAdapter.scala 111:25 chipyard.TestHarness.SmallBoomConfig.fir 394029:4]
  assign sim_serial_in_ready = rxfifo_io_enq_ready; // @[UARTAdapter.scala 119:26 chipyard.TestHarness.SmallBoomConfig.fir 394036:4]
  assign sim_serial_out_valid = txfifo_io_deq_valid; // @[UARTAdapter.scala 114:27 chipyard.TestHarness.SmallBoomConfig.fir 394032:4]
  assign sim_serial_out_bits = txfifo_io_deq_bits; // @[UARTAdapter.scala 113:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  always @(posedge clock) begin
    if (reset) begin // @[UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393878:4]
      txState <= 2'h0; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393878:4]
    end else if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.SmallBoomConfig.fir 393922:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.SmallBoomConfig.fir 393923:6]
        txState <= 2'h1; // @[UARTAdapter.scala 50:17 chipyard.TestHarness.SmallBoomConfig.fir 393925:8]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393930:6]
      if (txBaudWrap) begin // @[UARTAdapter.scala 54:24 chipyard.TestHarness.SmallBoomConfig.fir 393931:8]
        txState <= 2'h2; // @[UARTAdapter.scala 55:17 chipyard.TestHarness.SmallBoomConfig.fir 393932:10]
      end
    end else if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393937:8]
      txState <= _GEN_12;
    end else begin
      txState <= _GEN_14;
    end
    if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.SmallBoomConfig.fir 393922:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.SmallBoomConfig.fir 393923:6]
        txData <= 8'h0; // @[UARTAdapter.scala 49:17 chipyard.TestHarness.SmallBoomConfig.fir 393924:8]
      end
    end else if (!(_T_9)) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393930:6]
      if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393937:8]
        if (txfifo_io_enq_ready) begin // @[UARTAdapter.scala 59:34 chipyard.TestHarness.SmallBoomConfig.fir 393938:10]
          txData <= _txData_T_1; // @[UARTAdapter.scala 60:16 chipyard.TestHarness.SmallBoomConfig.fir 393941:12]
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393882:4]
      txDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393882:4]
    end else if (_T_1) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393885:4]
      txDataIdx <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393889:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393894:4]
      txBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393894:4]
    end else if (_T_3) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393897:4]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20 chipyard.TestHarness.SmallBoomConfig.fir 393902:6]
        txBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.SmallBoomConfig.fir 393903:8]
      end else begin
        txBaudCount <= _wrap_value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393901:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393911:4]
      txSlackCount <= 2'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393911:4]
    end else if (_T_7) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393914:4]
      txSlackCount <= _wrap_value_T_5; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393918:6]
    end
    if (reset) begin // @[UARTAdapter.scala 79:24 chipyard.TestHarness.SmallBoomConfig.fir 393964:4]
      rxState <= 2'h0; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.SmallBoomConfig.fir 393964:4]
    end else if (_T_17) begin // @[Conditional.scala 40:58 chipyard.TestHarness.SmallBoomConfig.fir 393993:4]
      if (_T_18) begin // @[UARTAdapter.scala 89:48 chipyard.TestHarness.SmallBoomConfig.fir 393996:6]
        rxState <= 2'h1; // @[UARTAdapter.scala 90:17 chipyard.TestHarness.SmallBoomConfig.fir 393997:8]
      end
    end else if (_T_19) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 394002:6]
      if (rxBaudWrap) begin // @[UARTAdapter.scala 95:24 chipyard.TestHarness.SmallBoomConfig.fir 394004:8]
        rxState <= 2'h2; // @[UARTAdapter.scala 96:17 chipyard.TestHarness.SmallBoomConfig.fir 394005:10]
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 394010:8]
      rxState <= _GEN_28;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393965:4]
      rxBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393965:4]
    end else if (txfifo_io_enq_ready) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393968:4]
      if (wrap_wrap_3) begin // @[Counter.scala 86:20 chipyard.TestHarness.SmallBoomConfig.fir 393973:6]
        rxBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.SmallBoomConfig.fir 393974:8]
      end else begin
        rxBaudCount <= _wrap_value_T_7; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393972:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393981:4]
      rxDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393981:4]
    end else if (_T_16) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393984:4]
      rxDataIdx <= _wrap_value_T_9; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393988:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  txState = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  txData = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  txDataIdx = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  txBaudCount = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  txSlackCount = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  rxState = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  rxBaudCount = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  rxDataIdx = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 394038:2]
  input   clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 394039:4]
  input   reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 394040:4]
  output  io_success // @[chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
);
  wire  chiptop_jtag_TCK; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_jtag_TMS; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_jtag_TDI; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_jtag_TDO_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_jtag_TDO_driven; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_serial_tl_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_serial_tl_bits_in_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_serial_tl_bits_in_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_serial_tl_bits_in_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_serial_tl_bits_out_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_serial_tl_bits_out_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_serial_tl_bits_out_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_reset; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_aw_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_aw_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [31:0] chiptop_axi4_mem_0_bits_aw_bits_addr; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [7:0] chiptop_axi4_mem_0_bits_aw_bits_len; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [2:0] chiptop_axi4_mem_0_bits_aw_bits_size; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [1:0] chiptop_axi4_mem_0_bits_aw_bits_burst; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_aw_bits_lock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_cache; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [2:0] chiptop_axi4_mem_0_bits_aw_bits_prot; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_qos; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_w_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_w_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [63:0] chiptop_axi4_mem_0_bits_w_bits_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [7:0] chiptop_axi4_mem_0_bits_w_bits_strb; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_w_bits_last; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_b_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_b_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_axi4_mem_0_bits_b_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [1:0] chiptop_axi4_mem_0_bits_b_bits_resp; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_ar_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_ar_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [31:0] chiptop_axi4_mem_0_bits_ar_bits_addr; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [7:0] chiptop_axi4_mem_0_bits_ar_bits_len; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [2:0] chiptop_axi4_mem_0_bits_ar_bits_size; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [1:0] chiptop_axi4_mem_0_bits_ar_bits_burst; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_ar_bits_lock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_cache; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [2:0] chiptop_axi4_mem_0_bits_ar_bits_prot; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_qos; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_r_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_r_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [3:0] chiptop_axi4_mem_0_bits_r_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [63:0] chiptop_axi4_mem_0_bits_r_bits_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire [1:0] chiptop_axi4_mem_0_bits_r_bits_resp; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_axi4_mem_0_bits_r_bits_last; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_uart_0_txd; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_uart_0_rxd; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_reset_wire_reset; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  chiptop_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
  wire  SimJTAG_clock; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_reset; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_jtag_TRSTn; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_jtag_TCK; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_jtag_TMS; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_jtag_TDI; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_jtag_TDO_data; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_jtag_TDO_driven; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_enable; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire  SimJTAG_init_done; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire [31:0] SimJTAG_exit; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 394072:4]
  wire  ram_clock; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_reset; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_io_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_io_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire [3:0] ram_io_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_io_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_io_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire [3:0] ram_io_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_io_tsi_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire [31:0] ram_io_tsi_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_io_tsi_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire [31:0] ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
  wire  success_sim_clock; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire  success_sim_reset; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire  success_sim_serial_in_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire  success_sim_serial_in_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire [31:0] success_sim_serial_in_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire  success_sim_serial_out_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire  success_sim_serial_out_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire [31:0] success_sim_serial_out_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire  success_sim_exit; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
  wire  simdram_clock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_reset; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_aw_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_aw_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [3:0] simdram_axi_aw_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [31:0] simdram_axi_aw_bits_addr; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [7:0] simdram_axi_aw_bits_len; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [2:0] simdram_axi_aw_bits_size; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [1:0] simdram_axi_aw_bits_burst; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_aw_bits_lock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [3:0] simdram_axi_aw_bits_cache; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [2:0] simdram_axi_aw_bits_prot; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [3:0] simdram_axi_aw_bits_qos; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_w_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_w_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [63:0] simdram_axi_w_bits_data; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [7:0] simdram_axi_w_bits_strb; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_w_bits_last; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_b_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_b_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [3:0] simdram_axi_b_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [1:0] simdram_axi_b_bits_resp; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_ar_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_ar_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [3:0] simdram_axi_ar_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [31:0] simdram_axi_ar_bits_addr; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [7:0] simdram_axi_ar_bits_len; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [2:0] simdram_axi_ar_bits_size; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [1:0] simdram_axi_ar_bits_burst; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_ar_bits_lock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [3:0] simdram_axi_ar_bits_cache; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [2:0] simdram_axi_ar_bits_prot; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [3:0] simdram_axi_ar_bits_qos; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_r_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_r_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [3:0] simdram_axi_r_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [63:0] simdram_axi_r_bits_data; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire [1:0] simdram_axi_r_bits_resp; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  simdram_axi_r_bits_last; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
  wire  uart_sim_0_clock; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394125:4]
  wire  uart_sim_0_reset; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394125:4]
  wire  uart_sim_0_io_uart_txd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394125:4]
  wire  uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394125:4]
  wire  dtm_success = SimJTAG_exit == 32'h1; // @[Periphery.scala 233:26 chipyard.TestHarness.SmallBoomConfig.fir 394076:4]
  wire  _T_2 = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.SmallBoomConfig.fir 394064:4]
  wire  _T_3 = SimJTAG_exit >= 32'h2; // @[Periphery.scala 234:19 chipyard.TestHarness.SmallBoomConfig.fir 394078:4]
  wire [31:0] _T_4 = {{1'd0}, SimJTAG_exit[31:1]}; // @[Periphery.scala 235:59 chipyard.TestHarness.SmallBoomConfig.fir 394080:6]
  ChipTop chiptop ( // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 394043:4]
    .jtag_TCK(chiptop_jtag_TCK),
    .jtag_TMS(chiptop_jtag_TMS),
    .jtag_TDI(chiptop_jtag_TDI),
    .jtag_TDO_data(chiptop_jtag_TDO_data),
    .jtag_TDO_driven(chiptop_jtag_TDO_driven),
    .serial_tl_clock(chiptop_serial_tl_clock),
    .serial_tl_bits_in_ready(chiptop_serial_tl_bits_in_ready),
    .serial_tl_bits_in_valid(chiptop_serial_tl_bits_in_valid),
    .serial_tl_bits_in_bits(chiptop_serial_tl_bits_in_bits),
    .serial_tl_bits_out_ready(chiptop_serial_tl_bits_out_ready),
    .serial_tl_bits_out_valid(chiptop_serial_tl_bits_out_valid),
    .serial_tl_bits_out_bits(chiptop_serial_tl_bits_out_bits),
    .axi4_mem_0_clock(chiptop_axi4_mem_0_clock),
    .axi4_mem_0_reset(chiptop_axi4_mem_0_reset),
    .axi4_mem_0_bits_aw_ready(chiptop_axi4_mem_0_bits_aw_ready),
    .axi4_mem_0_bits_aw_valid(chiptop_axi4_mem_0_bits_aw_valid),
    .axi4_mem_0_bits_aw_bits_id(chiptop_axi4_mem_0_bits_aw_bits_id),
    .axi4_mem_0_bits_aw_bits_addr(chiptop_axi4_mem_0_bits_aw_bits_addr),
    .axi4_mem_0_bits_aw_bits_len(chiptop_axi4_mem_0_bits_aw_bits_len),
    .axi4_mem_0_bits_aw_bits_size(chiptop_axi4_mem_0_bits_aw_bits_size),
    .axi4_mem_0_bits_aw_bits_burst(chiptop_axi4_mem_0_bits_aw_bits_burst),
    .axi4_mem_0_bits_aw_bits_lock(chiptop_axi4_mem_0_bits_aw_bits_lock),
    .axi4_mem_0_bits_aw_bits_cache(chiptop_axi4_mem_0_bits_aw_bits_cache),
    .axi4_mem_0_bits_aw_bits_prot(chiptop_axi4_mem_0_bits_aw_bits_prot),
    .axi4_mem_0_bits_aw_bits_qos(chiptop_axi4_mem_0_bits_aw_bits_qos),
    .axi4_mem_0_bits_w_ready(chiptop_axi4_mem_0_bits_w_ready),
    .axi4_mem_0_bits_w_valid(chiptop_axi4_mem_0_bits_w_valid),
    .axi4_mem_0_bits_w_bits_data(chiptop_axi4_mem_0_bits_w_bits_data),
    .axi4_mem_0_bits_w_bits_strb(chiptop_axi4_mem_0_bits_w_bits_strb),
    .axi4_mem_0_bits_w_bits_last(chiptop_axi4_mem_0_bits_w_bits_last),
    .axi4_mem_0_bits_b_ready(chiptop_axi4_mem_0_bits_b_ready),
    .axi4_mem_0_bits_b_valid(chiptop_axi4_mem_0_bits_b_valid),
    .axi4_mem_0_bits_b_bits_id(chiptop_axi4_mem_0_bits_b_bits_id),
    .axi4_mem_0_bits_b_bits_resp(chiptop_axi4_mem_0_bits_b_bits_resp),
    .axi4_mem_0_bits_ar_ready(chiptop_axi4_mem_0_bits_ar_ready),
    .axi4_mem_0_bits_ar_valid(chiptop_axi4_mem_0_bits_ar_valid),
    .axi4_mem_0_bits_ar_bits_id(chiptop_axi4_mem_0_bits_ar_bits_id),
    .axi4_mem_0_bits_ar_bits_addr(chiptop_axi4_mem_0_bits_ar_bits_addr),
    .axi4_mem_0_bits_ar_bits_len(chiptop_axi4_mem_0_bits_ar_bits_len),
    .axi4_mem_0_bits_ar_bits_size(chiptop_axi4_mem_0_bits_ar_bits_size),
    .axi4_mem_0_bits_ar_bits_burst(chiptop_axi4_mem_0_bits_ar_bits_burst),
    .axi4_mem_0_bits_ar_bits_lock(chiptop_axi4_mem_0_bits_ar_bits_lock),
    .axi4_mem_0_bits_ar_bits_cache(chiptop_axi4_mem_0_bits_ar_bits_cache),
    .axi4_mem_0_bits_ar_bits_prot(chiptop_axi4_mem_0_bits_ar_bits_prot),
    .axi4_mem_0_bits_ar_bits_qos(chiptop_axi4_mem_0_bits_ar_bits_qos),
    .axi4_mem_0_bits_r_ready(chiptop_axi4_mem_0_bits_r_ready),
    .axi4_mem_0_bits_r_valid(chiptop_axi4_mem_0_bits_r_valid),
    .axi4_mem_0_bits_r_bits_id(chiptop_axi4_mem_0_bits_r_bits_id),
    .axi4_mem_0_bits_r_bits_data(chiptop_axi4_mem_0_bits_r_bits_data),
    .axi4_mem_0_bits_r_bits_resp(chiptop_axi4_mem_0_bits_r_bits_resp),
    .axi4_mem_0_bits_r_bits_last(chiptop_axi4_mem_0_bits_r_bits_last),
    .uart_0_txd(chiptop_uart_0_txd),
    .uart_0_rxd(chiptop_uart_0_rxd),
    .reset_wire_reset(chiptop_reset_wire_reset),
    .clock(chiptop_clock)
  );
  SimJTAG #(.TICK_DELAY(3)) SimJTAG ( // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 394055:4]
    .clock(SimJTAG_clock),
    .reset(SimJTAG_reset),
    .jtag_TRSTn(SimJTAG_jtag_TRSTn),
    .jtag_TCK(SimJTAG_jtag_TCK),
    .jtag_TMS(SimJTAG_jtag_TMS),
    .jtag_TDI(SimJTAG_jtag_TDI),
    .jtag_TDO_data(SimJTAG_jtag_TDO_data),
    .jtag_TDO_driven(SimJTAG_jtag_TDO_driven),
    .enable(SimJTAG_enable),
    .init_done(SimJTAG_init_done),
    .exit(SimJTAG_exit)
  );
  plusarg_reader #(.FORMAT("jtag_rbb_enable=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 394072:4]
    .out(plusarg_reader_out)
  );
  SerialRAM_inTestHarness ram ( // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394092:4]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_ser_in_ready(ram_io_ser_in_ready),
    .io_ser_in_valid(ram_io_ser_in_valid),
    .io_ser_in_bits(ram_io_ser_in_bits),
    .io_ser_out_ready(ram_io_ser_out_ready),
    .io_ser_out_valid(ram_io_ser_out_valid),
    .io_ser_out_bits(ram_io_ser_out_bits),
    .io_tsi_ser_in_ready(ram_io_tsi_ser_in_ready),
    .io_tsi_ser_in_valid(ram_io_tsi_ser_in_valid),
    .io_tsi_ser_in_bits(ram_io_tsi_ser_in_bits),
    .io_tsi_ser_out_ready(ram_io_tsi_ser_out_ready),
    .io_tsi_ser_out_valid(ram_io_tsi_ser_out_valid),
    .io_tsi_ser_out_bits(ram_io_tsi_ser_out_bits)
  );
  SimSerial success_sim ( // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394102:4]
    .clock(success_sim_clock),
    .reset(success_sim_reset),
    .serial_in_ready(success_sim_serial_in_ready),
    .serial_in_valid(success_sim_serial_in_valid),
    .serial_in_bits(success_sim_serial_in_bits),
    .serial_out_ready(success_sim_serial_out_ready),
    .serial_out_valid(success_sim_serial_out_valid),
    .serial_out_bits(success_sim_serial_out_bits),
    .exit(success_sim_exit)
  );
  SimDRAM #(.LINE_SIZE(64), .ID_BITS(4), .ADDR_BITS(32), .MEM_SIZE(268435456), .DATA_BITS(64)) simdram ( // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394118:4]
    .clock(simdram_clock),
    .reset(simdram_reset),
    .axi_aw_ready(simdram_axi_aw_ready),
    .axi_aw_valid(simdram_axi_aw_valid),
    .axi_aw_bits_id(simdram_axi_aw_bits_id),
    .axi_aw_bits_addr(simdram_axi_aw_bits_addr),
    .axi_aw_bits_len(simdram_axi_aw_bits_len),
    .axi_aw_bits_size(simdram_axi_aw_bits_size),
    .axi_aw_bits_burst(simdram_axi_aw_bits_burst),
    .axi_aw_bits_lock(simdram_axi_aw_bits_lock),
    .axi_aw_bits_cache(simdram_axi_aw_bits_cache),
    .axi_aw_bits_prot(simdram_axi_aw_bits_prot),
    .axi_aw_bits_qos(simdram_axi_aw_bits_qos),
    .axi_w_ready(simdram_axi_w_ready),
    .axi_w_valid(simdram_axi_w_valid),
    .axi_w_bits_data(simdram_axi_w_bits_data),
    .axi_w_bits_strb(simdram_axi_w_bits_strb),
    .axi_w_bits_last(simdram_axi_w_bits_last),
    .axi_b_ready(simdram_axi_b_ready),
    .axi_b_valid(simdram_axi_b_valid),
    .axi_b_bits_id(simdram_axi_b_bits_id),
    .axi_b_bits_resp(simdram_axi_b_bits_resp),
    .axi_ar_ready(simdram_axi_ar_ready),
    .axi_ar_valid(simdram_axi_ar_valid),
    .axi_ar_bits_id(simdram_axi_ar_bits_id),
    .axi_ar_bits_addr(simdram_axi_ar_bits_addr),
    .axi_ar_bits_len(simdram_axi_ar_bits_len),
    .axi_ar_bits_size(simdram_axi_ar_bits_size),
    .axi_ar_bits_burst(simdram_axi_ar_bits_burst),
    .axi_ar_bits_lock(simdram_axi_ar_bits_lock),
    .axi_ar_bits_cache(simdram_axi_ar_bits_cache),
    .axi_ar_bits_prot(simdram_axi_ar_bits_prot),
    .axi_ar_bits_qos(simdram_axi_ar_bits_qos),
    .axi_r_ready(simdram_axi_r_ready),
    .axi_r_valid(simdram_axi_r_valid),
    .axi_r_bits_id(simdram_axi_r_bits_id),
    .axi_r_bits_data(simdram_axi_r_bits_data),
    .axi_r_bits_resp(simdram_axi_r_bits_resp),
    .axi_r_bits_last(simdram_axi_r_bits_last)
  );
  UARTAdapter_inTestHarness uart_sim_0 ( // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394125:4]
    .clock(uart_sim_0_clock),
    .reset(uart_sim_0_reset),
    .io_uart_txd(uart_sim_0_io_uart_txd),
    .io_uart_rxd(uart_sim_0_io_uart_rxd)
  );
  assign io_success = success_sim_exit | dtm_success; // @[HarnessBinders.scala 236:22 chipyard.TestHarness.SmallBoomConfig.fir 394115:4 HarnessBinders.scala 236:35 chipyard.TestHarness.SmallBoomConfig.fir 394116:6]
  assign chiptop_jtag_TCK = SimJTAG_jtag_TCK; // @[Periphery.scala 220:15 chipyard.TestHarness.SmallBoomConfig.fir 394065:4]
  assign chiptop_jtag_TMS = SimJTAG_jtag_TMS; // @[Periphery.scala 221:15 chipyard.TestHarness.SmallBoomConfig.fir 394066:4]
  assign chiptop_jtag_TDI = SimJTAG_jtag_TDI; // @[Periphery.scala 222:15 chipyard.TestHarness.SmallBoomConfig.fir 394067:4]
  assign chiptop_serial_tl_bits_in_valid = ram_io_ser_in_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394099:4]
  assign chiptop_serial_tl_bits_in_bits = ram_io_ser_in_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394098:4]
  assign chiptop_serial_tl_bits_out_ready = ram_io_ser_out_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394097:4]
  assign chiptop_axi4_mem_0_bits_aw_ready = simdram_axi_aw_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_w_ready = simdram_axi_w_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_b_valid = simdram_axi_b_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_b_bits_id = simdram_axi_b_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_b_bits_resp = simdram_axi_b_bits_resp; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_ar_ready = simdram_axi_ar_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_r_valid = simdram_axi_r_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_r_bits_id = simdram_axi_r_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_r_bits_data = simdram_axi_r_bits_data; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_r_bits_resp = simdram_axi_r_bits_resp; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_axi4_mem_0_bits_r_bits_last = simdram_axi_r_bits_last; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign chiptop_uart_0_rxd = uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 135:18 chipyard.TestHarness.SmallBoomConfig.fir 394129:4]
  assign chiptop_reset_wire_reset = reset; // @[TestHarness.scala 41:24 chipyard.TestHarness.SmallBoomConfig.fir 394047:4]
  assign chiptop_clock = clock; // @[Clocks.scala 106:18 chipyard.TestHarness.SmallBoomConfig.fir 394049:4]
  assign SimJTAG_clock = clock; // @[Periphery.scala 225:14 chipyard.TestHarness.SmallBoomConfig.fir 394070:4]
  assign SimJTAG_reset = reset; // @[HarnessBinders.scala 190:97 chipyard.TestHarness.SmallBoomConfig.fir 394062:4]
  assign SimJTAG_jtag_TDO_data = chiptop_jtag_TDO_data; // @[Periphery.scala 223:17 chipyard.TestHarness.SmallBoomConfig.fir 394069:4]
  assign SimJTAG_jtag_TDO_driven = chiptop_jtag_TDO_driven; // @[Periphery.scala 223:17 chipyard.TestHarness.SmallBoomConfig.fir 394068:4]
  assign SimJTAG_enable = plusarg_reader_out[0]; // @[Periphery.scala 228:18 chipyard.TestHarness.SmallBoomConfig.fir 394074:4]
  assign SimJTAG_init_done = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.SmallBoomConfig.fir 394064:4]
  assign ram_clock = chiptop_serial_tl_clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 394093:4]
  assign ram_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 394045:4 chipyard.TestHarness.SmallBoomConfig.fir 394046:4]
  assign ram_io_ser_in_ready = chiptop_serial_tl_bits_in_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394100:4]
  assign ram_io_ser_out_valid = chiptop_serial_tl_bits_out_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394096:4]
  assign ram_io_ser_out_bits = chiptop_serial_tl_bits_out_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394095:4]
  assign ram_io_tsi_ser_in_valid = success_sim_serial_in_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394113:4]
  assign ram_io_tsi_ser_in_bits = success_sim_serial_in_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394112:4]
  assign ram_io_tsi_ser_out_ready = success_sim_serial_out_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394111:4]
  assign success_sim_clock = chiptop_serial_tl_clock; // @[SerialAdapter.scala 38:20 chipyard.TestHarness.SmallBoomConfig.fir 394107:4]
  assign success_sim_reset = reset; // @[HarnessBinders.scala 235:103 chipyard.TestHarness.SmallBoomConfig.fir 394101:4]
  assign success_sim_serial_in_ready = ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394114:4]
  assign success_sim_serial_out_valid = ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394110:4]
  assign success_sim_serial_out_bits = ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394109:4]
  assign simdram_clock = chiptop_axi4_mem_0_clock; // @[HarnessBinders.scala 148:20 chipyard.TestHarness.SmallBoomConfig.fir 394123:4]
  assign simdram_reset = chiptop_axi4_mem_0_reset; // @[HarnessBinders.scala 149:20 chipyard.TestHarness.SmallBoomConfig.fir 394124:4]
  assign simdram_axi_aw_valid = chiptop_axi4_mem_0_bits_aw_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_id = chiptop_axi4_mem_0_bits_aw_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_addr = chiptop_axi4_mem_0_bits_aw_bits_addr; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_len = chiptop_axi4_mem_0_bits_aw_bits_len; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_size = chiptop_axi4_mem_0_bits_aw_bits_size; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_burst = chiptop_axi4_mem_0_bits_aw_bits_burst; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_lock = chiptop_axi4_mem_0_bits_aw_bits_lock; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_cache = chiptop_axi4_mem_0_bits_aw_bits_cache; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_prot = chiptop_axi4_mem_0_bits_aw_bits_prot; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_aw_bits_qos = chiptop_axi4_mem_0_bits_aw_bits_qos; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_w_valid = chiptop_axi4_mem_0_bits_w_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_w_bits_data = chiptop_axi4_mem_0_bits_w_bits_data; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_w_bits_strb = chiptop_axi4_mem_0_bits_w_bits_strb; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_w_bits_last = chiptop_axi4_mem_0_bits_w_bits_last; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_b_ready = chiptop_axi4_mem_0_bits_b_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_valid = chiptop_axi4_mem_0_bits_ar_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_id = chiptop_axi4_mem_0_bits_ar_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_addr = chiptop_axi4_mem_0_bits_ar_bits_addr; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_len = chiptop_axi4_mem_0_bits_ar_bits_len; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_size = chiptop_axi4_mem_0_bits_ar_bits_size; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_burst = chiptop_axi4_mem_0_bits_ar_bits_burst; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_lock = chiptop_axi4_mem_0_bits_ar_bits_lock; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_cache = chiptop_axi4_mem_0_bits_ar_bits_cache; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_prot = chiptop_axi4_mem_0_bits_ar_bits_prot; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_ar_bits_qos = chiptop_axi4_mem_0_bits_ar_bits_qos; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign simdram_axi_r_ready = chiptop_axi4_mem_0_bits_r_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394122:4]
  assign uart_sim_0_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 394126:4]
  assign uart_sim_0_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 394127:4]
  assign uart_sim_0_io_uart_txd = chiptop_uart_0_txd; // @[UARTAdapter.scala 134:28 chipyard.TestHarness.SmallBoomConfig.fir 394128:4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fwrite(32'h80000002,"*** FAILED *** (exit code = %d)\n",_T_4); // @[Periphery.scala 235:13 chipyard.TestHarness.SmallBoomConfig.fir 394084:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fatal; // @[Periphery.scala 236:11 chipyard.TestHarness.SmallBoomConfig.fir 394089:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module mem_inTestHarness(
  input  [8:0] RW0_addr,
  input        RW0_en,
  input        RW0_clk,
  input        RW0_wmode,
  input  [7:0] RW0_wdata_0,
  input  [7:0] RW0_wdata_1,
  input  [7:0] RW0_wdata_2,
  input  [7:0] RW0_wdata_3,
  input  [7:0] RW0_wdata_4,
  input  [7:0] RW0_wdata_5,
  input  [7:0] RW0_wdata_6,
  input  [7:0] RW0_wdata_7,
  output [7:0] RW0_rdata_0,
  output [7:0] RW0_rdata_1,
  output [7:0] RW0_rdata_2,
  output [7:0] RW0_rdata_3,
  output [7:0] RW0_rdata_4,
  output [7:0] RW0_rdata_5,
  output [7:0] RW0_rdata_6,
  output [7:0] RW0_rdata_7,
  input        RW0_wmask_0,
  input        RW0_wmask_1,
  input        RW0_wmask_2,
  input        RW0_wmask_3,
  input        RW0_wmask_4,
  input        RW0_wmask_5,
  input        RW0_wmask_6,
  input        RW0_wmask_7
);
  wire [8:0] mem_ext_RW0_addr;
  wire  mem_ext_RW0_en;
  wire  mem_ext_RW0_clk;
  wire  mem_ext_RW0_wmode;
  wire [63:0] mem_ext_RW0_wdata;
  wire [63:0] mem_ext_RW0_rdata;
  wire [7:0] mem_ext_RW0_wmask;
  wire [31:0] _GEN_4 = {RW0_wdata_7,RW0_wdata_6,RW0_wdata_5,RW0_wdata_4};
  wire [31:0] _GEN_5 = {RW0_wdata_3,RW0_wdata_2,RW0_wdata_1,RW0_wdata_0};
  wire [3:0] _GEN_10 = {RW0_wmask_7,RW0_wmask_6,RW0_wmask_5,RW0_wmask_4};
  wire [3:0] _GEN_11 = {RW0_wmask_3,RW0_wmask_2,RW0_wmask_1,RW0_wmask_0};
  mem_ext mem_ext (
    .RW0_addr(mem_ext_RW0_addr),
    .RW0_en(mem_ext_RW0_en),
    .RW0_clk(mem_ext_RW0_clk),
    .RW0_wmode(mem_ext_RW0_wmode),
    .RW0_wdata(mem_ext_RW0_wdata),
    .RW0_rdata(mem_ext_RW0_rdata),
    .RW0_wmask(mem_ext_RW0_wmask)
  );
  assign mem_ext_RW0_clk = RW0_clk;
  assign mem_ext_RW0_en = RW0_en;
  assign mem_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = mem_ext_RW0_rdata[7:0];
  assign RW0_rdata_1 = mem_ext_RW0_rdata[15:8];
  assign RW0_rdata_2 = mem_ext_RW0_rdata[23:16];
  assign RW0_rdata_3 = mem_ext_RW0_rdata[31:24];
  assign RW0_rdata_4 = mem_ext_RW0_rdata[39:32];
  assign RW0_rdata_5 = mem_ext_RW0_rdata[47:40];
  assign RW0_rdata_6 = mem_ext_RW0_rdata[55:48];
  assign RW0_rdata_7 = mem_ext_RW0_rdata[63:56];
  assign mem_ext_RW0_wmode = RW0_wmode;
  assign mem_ext_RW0_wdata = {_GEN_4,_GEN_5};
  assign mem_ext_RW0_wmask = {_GEN_10,_GEN_11};
endmodule
